module rom_go (clock, address, q);
input clock;
output [0:0] q;
input [15:0] address;
reg [0:0] dout;
reg [0:0] ram [65535:0];
assign q = dout;

initial begin
  ram[0]  = 1;
  ram[1]  = 1;
  ram[2]  = 1;
  ram[3]  = 1;
  ram[4]  = 1;
  ram[5]  = 1;
  ram[6]  = 1;
  ram[7]  = 1;
  ram[8]  = 1;
  ram[9]  = 1;
  ram[10]  = 1;
  ram[11]  = 1;
  ram[12]  = 1;
  ram[13]  = 1;
  ram[14]  = 1;
  ram[15]  = 1;
  ram[16]  = 1;
  ram[17]  = 1;
  ram[18]  = 1;
  ram[19]  = 1;
  ram[20]  = 1;
  ram[21]  = 1;
  ram[22]  = 1;
  ram[23]  = 1;
  ram[24]  = 1;
  ram[25]  = 1;
  ram[26]  = 1;
  ram[27]  = 1;
  ram[28]  = 1;
  ram[29]  = 1;
  ram[30]  = 1;
  ram[31]  = 1;
  ram[32]  = 1;
  ram[33]  = 1;
  ram[34]  = 1;
  ram[35]  = 1;
  ram[36]  = 1;
  ram[37]  = 1;
  ram[38]  = 1;
  ram[39]  = 1;
  ram[40]  = 1;
  ram[41]  = 1;
  ram[42]  = 1;
  ram[43]  = 1;
  ram[44]  = 1;
  ram[45]  = 1;
  ram[46]  = 1;
  ram[47]  = 1;
  ram[48]  = 1;
  ram[49]  = 1;
  ram[50]  = 1;
  ram[51]  = 1;
  ram[52]  = 1;
  ram[53]  = 1;
  ram[54]  = 1;
  ram[55]  = 1;
  ram[56]  = 1;
  ram[57]  = 1;
  ram[58]  = 1;
  ram[59]  = 1;
  ram[60]  = 1;
  ram[61]  = 1;
  ram[62]  = 1;
  ram[63]  = 1;
  ram[64]  = 1;
  ram[65]  = 1;
  ram[66]  = 1;
  ram[67]  = 1;
  ram[68]  = 1;
  ram[69]  = 1;
  ram[70]  = 1;
  ram[71]  = 1;
  ram[72]  = 1;
  ram[73]  = 1;
  ram[74]  = 1;
  ram[75]  = 1;
  ram[76]  = 1;
  ram[77]  = 1;
  ram[78]  = 1;
  ram[79]  = 1;
  ram[80]  = 1;
  ram[81]  = 1;
  ram[82]  = 1;
  ram[83]  = 1;
  ram[84]  = 1;
  ram[85]  = 1;
  ram[86]  = 1;
  ram[87]  = 1;
  ram[88]  = 1;
  ram[89]  = 1;
  ram[90]  = 1;
  ram[91]  = 1;
  ram[92]  = 1;
  ram[93]  = 1;
  ram[94]  = 1;
  ram[95]  = 1;
  ram[96]  = 1;
  ram[97]  = 1;
  ram[98]  = 1;
  ram[99]  = 1;
  ram[100]  = 1;
  ram[101]  = 1;
  ram[102]  = 1;
  ram[103]  = 1;
  ram[104]  = 1;
  ram[105]  = 1;
  ram[106]  = 1;
  ram[107]  = 1;
  ram[108]  = 1;
  ram[109]  = 1;
  ram[110]  = 1;
  ram[111]  = 1;
  ram[112]  = 1;
  ram[113]  = 1;
  ram[114]  = 1;
  ram[115]  = 1;
  ram[116]  = 1;
  ram[117]  = 1;
  ram[118]  = 1;
  ram[119]  = 1;
  ram[120]  = 1;
  ram[121]  = 1;
  ram[122]  = 1;
  ram[123]  = 1;
  ram[124]  = 1;
  ram[125]  = 1;
  ram[126]  = 1;
  ram[127]  = 1;
  ram[128]  = 1;
  ram[129]  = 1;
  ram[130]  = 1;
  ram[131]  = 1;
  ram[132]  = 1;
  ram[133]  = 1;
  ram[134]  = 1;
  ram[135]  = 1;
  ram[136]  = 1;
  ram[137]  = 1;
  ram[138]  = 1;
  ram[139]  = 1;
  ram[140]  = 1;
  ram[141]  = 1;
  ram[142]  = 1;
  ram[143]  = 1;
  ram[144]  = 1;
  ram[145]  = 1;
  ram[146]  = 1;
  ram[147]  = 1;
  ram[148]  = 1;
  ram[149]  = 1;
  ram[150]  = 1;
  ram[151]  = 1;
  ram[152]  = 1;
  ram[153]  = 1;
  ram[154]  = 1;
  ram[155]  = 1;
  ram[156]  = 1;
  ram[157]  = 1;
  ram[158]  = 1;
  ram[159]  = 1;
  ram[160]  = 1;
  ram[161]  = 1;
  ram[162]  = 1;
  ram[163]  = 1;
  ram[164]  = 1;
  ram[165]  = 1;
  ram[166]  = 1;
  ram[167]  = 1;
  ram[168]  = 1;
  ram[169]  = 1;
  ram[170]  = 1;
  ram[171]  = 1;
  ram[172]  = 1;
  ram[173]  = 1;
  ram[174]  = 1;
  ram[175]  = 1;
  ram[176]  = 1;
  ram[177]  = 1;
  ram[178]  = 1;
  ram[179]  = 1;
  ram[180]  = 1;
  ram[181]  = 1;
  ram[182]  = 1;
  ram[183]  = 1;
  ram[184]  = 1;
  ram[185]  = 1;
  ram[186]  = 1;
  ram[187]  = 1;
  ram[188]  = 1;
  ram[189]  = 1;
  ram[190]  = 1;
  ram[191]  = 1;
  ram[192]  = 1;
  ram[193]  = 1;
  ram[194]  = 1;
  ram[195]  = 1;
  ram[196]  = 1;
  ram[197]  = 1;
  ram[198]  = 1;
  ram[199]  = 1;
  ram[200]  = 1;
  ram[201]  = 1;
  ram[202]  = 1;
  ram[203]  = 1;
  ram[204]  = 1;
  ram[205]  = 1;
  ram[206]  = 1;
  ram[207]  = 1;
  ram[208]  = 1;
  ram[209]  = 1;
  ram[210]  = 1;
  ram[211]  = 1;
  ram[212]  = 1;
  ram[213]  = 1;
  ram[214]  = 1;
  ram[215]  = 1;
  ram[216]  = 1;
  ram[217]  = 1;
  ram[218]  = 1;
  ram[219]  = 1;
  ram[220]  = 1;
  ram[221]  = 1;
  ram[222]  = 1;
  ram[223]  = 1;
  ram[224]  = 1;
  ram[225]  = 1;
  ram[226]  = 1;
  ram[227]  = 1;
  ram[228]  = 1;
  ram[229]  = 1;
  ram[230]  = 1;
  ram[231]  = 1;
  ram[232]  = 1;
  ram[233]  = 1;
  ram[234]  = 1;
  ram[235]  = 1;
  ram[236]  = 1;
  ram[237]  = 1;
  ram[238]  = 1;
  ram[239]  = 1;
  ram[240]  = 1;
  ram[241]  = 1;
  ram[242]  = 1;
  ram[243]  = 1;
  ram[244]  = 1;
  ram[245]  = 1;
  ram[246]  = 1;
  ram[247]  = 1;
  ram[248]  = 1;
  ram[249]  = 1;
  ram[250]  = 1;
  ram[251]  = 1;
  ram[252]  = 1;
  ram[253]  = 1;
  ram[254]  = 1;
  ram[255]  = 1;
  ram[256]  = 1;
  ram[257]  = 1;
  ram[258]  = 1;
  ram[259]  = 1;
  ram[260]  = 1;
  ram[261]  = 1;
  ram[262]  = 1;
  ram[263]  = 1;
  ram[264]  = 1;
  ram[265]  = 1;
  ram[266]  = 1;
  ram[267]  = 1;
  ram[268]  = 1;
  ram[269]  = 1;
  ram[270]  = 1;
  ram[271]  = 1;
  ram[272]  = 1;
  ram[273]  = 1;
  ram[274]  = 1;
  ram[275]  = 1;
  ram[276]  = 1;
  ram[277]  = 1;
  ram[278]  = 1;
  ram[279]  = 1;
  ram[280]  = 1;
  ram[281]  = 1;
  ram[282]  = 1;
  ram[283]  = 1;
  ram[284]  = 1;
  ram[285]  = 1;
  ram[286]  = 1;
  ram[287]  = 1;
  ram[288]  = 1;
  ram[289]  = 1;
  ram[290]  = 1;
  ram[291]  = 1;
  ram[292]  = 1;
  ram[293]  = 1;
  ram[294]  = 1;
  ram[295]  = 1;
  ram[296]  = 1;
  ram[297]  = 1;
  ram[298]  = 1;
  ram[299]  = 1;
  ram[300]  = 1;
  ram[301]  = 1;
  ram[302]  = 1;
  ram[303]  = 1;
  ram[304]  = 1;
  ram[305]  = 1;
  ram[306]  = 1;
  ram[307]  = 1;
  ram[308]  = 1;
  ram[309]  = 1;
  ram[310]  = 1;
  ram[311]  = 1;
  ram[312]  = 1;
  ram[313]  = 1;
  ram[314]  = 1;
  ram[315]  = 1;
  ram[316]  = 1;
  ram[317]  = 1;
  ram[318]  = 1;
  ram[319]  = 1;
  ram[320]  = 1;
  ram[321]  = 1;
  ram[322]  = 1;
  ram[323]  = 1;
  ram[324]  = 1;
  ram[325]  = 1;
  ram[326]  = 1;
  ram[327]  = 1;
  ram[328]  = 1;
  ram[329]  = 1;
  ram[330]  = 1;
  ram[331]  = 1;
  ram[332]  = 1;
  ram[333]  = 1;
  ram[334]  = 1;
  ram[335]  = 1;
  ram[336]  = 1;
  ram[337]  = 1;
  ram[338]  = 1;
  ram[339]  = 1;
  ram[340]  = 1;
  ram[341]  = 1;
  ram[342]  = 1;
  ram[343]  = 1;
  ram[344]  = 1;
  ram[345]  = 1;
  ram[346]  = 1;
  ram[347]  = 1;
  ram[348]  = 1;
  ram[349]  = 1;
  ram[350]  = 1;
  ram[351]  = 1;
  ram[352]  = 1;
  ram[353]  = 1;
  ram[354]  = 1;
  ram[355]  = 1;
  ram[356]  = 1;
  ram[357]  = 1;
  ram[358]  = 1;
  ram[359]  = 1;
  ram[360]  = 1;
  ram[361]  = 1;
  ram[362]  = 1;
  ram[363]  = 1;
  ram[364]  = 1;
  ram[365]  = 1;
  ram[366]  = 1;
  ram[367]  = 1;
  ram[368]  = 1;
  ram[369]  = 1;
  ram[370]  = 1;
  ram[371]  = 1;
  ram[372]  = 1;
  ram[373]  = 1;
  ram[374]  = 1;
  ram[375]  = 1;
  ram[376]  = 1;
  ram[377]  = 1;
  ram[378]  = 1;
  ram[379]  = 1;
  ram[380]  = 1;
  ram[381]  = 1;
  ram[382]  = 1;
  ram[383]  = 1;
  ram[384]  = 1;
  ram[385]  = 1;
  ram[386]  = 1;
  ram[387]  = 1;
  ram[388]  = 1;
  ram[389]  = 1;
  ram[390]  = 1;
  ram[391]  = 1;
  ram[392]  = 1;
  ram[393]  = 1;
  ram[394]  = 1;
  ram[395]  = 1;
  ram[396]  = 1;
  ram[397]  = 1;
  ram[398]  = 1;
  ram[399]  = 1;
  ram[400]  = 1;
  ram[401]  = 1;
  ram[402]  = 1;
  ram[403]  = 1;
  ram[404]  = 1;
  ram[405]  = 1;
  ram[406]  = 1;
  ram[407]  = 1;
  ram[408]  = 1;
  ram[409]  = 1;
  ram[410]  = 1;
  ram[411]  = 1;
  ram[412]  = 1;
  ram[413]  = 1;
  ram[414]  = 1;
  ram[415]  = 1;
  ram[416]  = 1;
  ram[417]  = 1;
  ram[418]  = 1;
  ram[419]  = 1;
  ram[420]  = 1;
  ram[421]  = 1;
  ram[422]  = 1;
  ram[423]  = 1;
  ram[424]  = 1;
  ram[425]  = 1;
  ram[426]  = 1;
  ram[427]  = 1;
  ram[428]  = 1;
  ram[429]  = 1;
  ram[430]  = 1;
  ram[431]  = 1;
  ram[432]  = 1;
  ram[433]  = 1;
  ram[434]  = 1;
  ram[435]  = 1;
  ram[436]  = 1;
  ram[437]  = 1;
  ram[438]  = 1;
  ram[439]  = 1;
  ram[440]  = 1;
  ram[441]  = 1;
  ram[442]  = 1;
  ram[443]  = 1;
  ram[444]  = 1;
  ram[445]  = 1;
  ram[446]  = 1;
  ram[447]  = 1;
  ram[448]  = 1;
  ram[449]  = 1;
  ram[450]  = 1;
  ram[451]  = 1;
  ram[452]  = 1;
  ram[453]  = 1;
  ram[454]  = 1;
  ram[455]  = 1;
  ram[456]  = 1;
  ram[457]  = 1;
  ram[458]  = 1;
  ram[459]  = 1;
  ram[460]  = 1;
  ram[461]  = 1;
  ram[462]  = 1;
  ram[463]  = 1;
  ram[464]  = 1;
  ram[465]  = 1;
  ram[466]  = 1;
  ram[467]  = 1;
  ram[468]  = 1;
  ram[469]  = 1;
  ram[470]  = 1;
  ram[471]  = 1;
  ram[472]  = 1;
  ram[473]  = 1;
  ram[474]  = 1;
  ram[475]  = 1;
  ram[476]  = 1;
  ram[477]  = 1;
  ram[478]  = 1;
  ram[479]  = 1;
  ram[480]  = 1;
  ram[481]  = 1;
  ram[482]  = 1;
  ram[483]  = 1;
  ram[484]  = 1;
  ram[485]  = 1;
  ram[486]  = 1;
  ram[487]  = 1;
  ram[488]  = 1;
  ram[489]  = 1;
  ram[490]  = 1;
  ram[491]  = 1;
  ram[492]  = 1;
  ram[493]  = 1;
  ram[494]  = 1;
  ram[495]  = 1;
  ram[496]  = 1;
  ram[497]  = 1;
  ram[498]  = 1;
  ram[499]  = 1;
  ram[500]  = 1;
  ram[501]  = 1;
  ram[502]  = 1;
  ram[503]  = 1;
  ram[504]  = 1;
  ram[505]  = 1;
  ram[506]  = 1;
  ram[507]  = 1;
  ram[508]  = 1;
  ram[509]  = 1;
  ram[510]  = 1;
  ram[511]  = 1;
  ram[512]  = 1;
  ram[513]  = 1;
  ram[514]  = 1;
  ram[515]  = 1;
  ram[516]  = 1;
  ram[517]  = 1;
  ram[518]  = 1;
  ram[519]  = 1;
  ram[520]  = 1;
  ram[521]  = 1;
  ram[522]  = 1;
  ram[523]  = 1;
  ram[524]  = 1;
  ram[525]  = 1;
  ram[526]  = 1;
  ram[527]  = 1;
  ram[528]  = 1;
  ram[529]  = 1;
  ram[530]  = 1;
  ram[531]  = 1;
  ram[532]  = 1;
  ram[533]  = 1;
  ram[534]  = 1;
  ram[535]  = 1;
  ram[536]  = 1;
  ram[537]  = 1;
  ram[538]  = 1;
  ram[539]  = 1;
  ram[540]  = 1;
  ram[541]  = 1;
  ram[542]  = 1;
  ram[543]  = 1;
  ram[544]  = 1;
  ram[545]  = 1;
  ram[546]  = 1;
  ram[547]  = 1;
  ram[548]  = 1;
  ram[549]  = 1;
  ram[550]  = 1;
  ram[551]  = 1;
  ram[552]  = 1;
  ram[553]  = 1;
  ram[554]  = 1;
  ram[555]  = 1;
  ram[556]  = 1;
  ram[557]  = 1;
  ram[558]  = 1;
  ram[559]  = 1;
  ram[560]  = 1;
  ram[561]  = 1;
  ram[562]  = 1;
  ram[563]  = 1;
  ram[564]  = 1;
  ram[565]  = 1;
  ram[566]  = 1;
  ram[567]  = 1;
  ram[568]  = 1;
  ram[569]  = 1;
  ram[570]  = 1;
  ram[571]  = 1;
  ram[572]  = 1;
  ram[573]  = 1;
  ram[574]  = 1;
  ram[575]  = 1;
  ram[576]  = 1;
  ram[577]  = 1;
  ram[578]  = 1;
  ram[579]  = 1;
  ram[580]  = 1;
  ram[581]  = 1;
  ram[582]  = 1;
  ram[583]  = 1;
  ram[584]  = 1;
  ram[585]  = 1;
  ram[586]  = 1;
  ram[587]  = 1;
  ram[588]  = 1;
  ram[589]  = 1;
  ram[590]  = 1;
  ram[591]  = 1;
  ram[592]  = 1;
  ram[593]  = 1;
  ram[594]  = 1;
  ram[595]  = 1;
  ram[596]  = 1;
  ram[597]  = 1;
  ram[598]  = 1;
  ram[599]  = 1;
  ram[600]  = 1;
  ram[601]  = 1;
  ram[602]  = 1;
  ram[603]  = 1;
  ram[604]  = 1;
  ram[605]  = 1;
  ram[606]  = 1;
  ram[607]  = 1;
  ram[608]  = 1;
  ram[609]  = 1;
  ram[610]  = 1;
  ram[611]  = 1;
  ram[612]  = 1;
  ram[613]  = 1;
  ram[614]  = 1;
  ram[615]  = 1;
  ram[616]  = 1;
  ram[617]  = 1;
  ram[618]  = 1;
  ram[619]  = 1;
  ram[620]  = 1;
  ram[621]  = 1;
  ram[622]  = 1;
  ram[623]  = 1;
  ram[624]  = 1;
  ram[625]  = 1;
  ram[626]  = 1;
  ram[627]  = 1;
  ram[628]  = 1;
  ram[629]  = 1;
  ram[630]  = 1;
  ram[631]  = 1;
  ram[632]  = 1;
  ram[633]  = 1;
  ram[634]  = 1;
  ram[635]  = 1;
  ram[636]  = 1;
  ram[637]  = 1;
  ram[638]  = 1;
  ram[639]  = 1;
  ram[640]  = 1;
  ram[641]  = 1;
  ram[642]  = 1;
  ram[643]  = 1;
  ram[644]  = 1;
  ram[645]  = 1;
  ram[646]  = 1;
  ram[647]  = 1;
  ram[648]  = 1;
  ram[649]  = 1;
  ram[650]  = 1;
  ram[651]  = 1;
  ram[652]  = 1;
  ram[653]  = 1;
  ram[654]  = 1;
  ram[655]  = 1;
  ram[656]  = 1;
  ram[657]  = 1;
  ram[658]  = 1;
  ram[659]  = 1;
  ram[660]  = 1;
  ram[661]  = 1;
  ram[662]  = 1;
  ram[663]  = 1;
  ram[664]  = 1;
  ram[665]  = 1;
  ram[666]  = 1;
  ram[667]  = 1;
  ram[668]  = 1;
  ram[669]  = 1;
  ram[670]  = 1;
  ram[671]  = 1;
  ram[672]  = 1;
  ram[673]  = 1;
  ram[674]  = 1;
  ram[675]  = 1;
  ram[676]  = 1;
  ram[677]  = 1;
  ram[678]  = 1;
  ram[679]  = 1;
  ram[680]  = 1;
  ram[681]  = 1;
  ram[682]  = 1;
  ram[683]  = 1;
  ram[684]  = 1;
  ram[685]  = 1;
  ram[686]  = 1;
  ram[687]  = 1;
  ram[688]  = 1;
  ram[689]  = 1;
  ram[690]  = 1;
  ram[691]  = 1;
  ram[692]  = 1;
  ram[693]  = 1;
  ram[694]  = 1;
  ram[695]  = 1;
  ram[696]  = 1;
  ram[697]  = 1;
  ram[698]  = 1;
  ram[699]  = 1;
  ram[700]  = 1;
  ram[701]  = 1;
  ram[702]  = 1;
  ram[703]  = 1;
  ram[704]  = 1;
  ram[705]  = 1;
  ram[706]  = 1;
  ram[707]  = 1;
  ram[708]  = 1;
  ram[709]  = 1;
  ram[710]  = 1;
  ram[711]  = 1;
  ram[712]  = 1;
  ram[713]  = 1;
  ram[714]  = 1;
  ram[715]  = 1;
  ram[716]  = 1;
  ram[717]  = 1;
  ram[718]  = 1;
  ram[719]  = 1;
  ram[720]  = 1;
  ram[721]  = 1;
  ram[722]  = 1;
  ram[723]  = 1;
  ram[724]  = 1;
  ram[725]  = 1;
  ram[726]  = 1;
  ram[727]  = 1;
  ram[728]  = 1;
  ram[729]  = 1;
  ram[730]  = 1;
  ram[731]  = 1;
  ram[732]  = 1;
  ram[733]  = 1;
  ram[734]  = 1;
  ram[735]  = 1;
  ram[736]  = 1;
  ram[737]  = 1;
  ram[738]  = 1;
  ram[739]  = 1;
  ram[740]  = 1;
  ram[741]  = 1;
  ram[742]  = 1;
  ram[743]  = 1;
  ram[744]  = 1;
  ram[745]  = 1;
  ram[746]  = 1;
  ram[747]  = 1;
  ram[748]  = 1;
  ram[749]  = 1;
  ram[750]  = 1;
  ram[751]  = 1;
  ram[752]  = 1;
  ram[753]  = 1;
  ram[754]  = 1;
  ram[755]  = 1;
  ram[756]  = 1;
  ram[757]  = 1;
  ram[758]  = 1;
  ram[759]  = 1;
  ram[760]  = 1;
  ram[761]  = 1;
  ram[762]  = 1;
  ram[763]  = 1;
  ram[764]  = 1;
  ram[765]  = 1;
  ram[766]  = 1;
  ram[767]  = 1;
  ram[768]  = 1;
  ram[769]  = 1;
  ram[770]  = 1;
  ram[771]  = 1;
  ram[772]  = 1;
  ram[773]  = 1;
  ram[774]  = 1;
  ram[775]  = 1;
  ram[776]  = 1;
  ram[777]  = 1;
  ram[778]  = 1;
  ram[779]  = 1;
  ram[780]  = 1;
  ram[781]  = 1;
  ram[782]  = 1;
  ram[783]  = 1;
  ram[784]  = 1;
  ram[785]  = 1;
  ram[786]  = 1;
  ram[787]  = 1;
  ram[788]  = 1;
  ram[789]  = 1;
  ram[790]  = 1;
  ram[791]  = 1;
  ram[792]  = 1;
  ram[793]  = 1;
  ram[794]  = 1;
  ram[795]  = 1;
  ram[796]  = 1;
  ram[797]  = 1;
  ram[798]  = 1;
  ram[799]  = 1;
  ram[800]  = 1;
  ram[801]  = 1;
  ram[802]  = 1;
  ram[803]  = 1;
  ram[804]  = 1;
  ram[805]  = 1;
  ram[806]  = 1;
  ram[807]  = 1;
  ram[808]  = 1;
  ram[809]  = 1;
  ram[810]  = 1;
  ram[811]  = 1;
  ram[812]  = 1;
  ram[813]  = 1;
  ram[814]  = 1;
  ram[815]  = 1;
  ram[816]  = 1;
  ram[817]  = 1;
  ram[818]  = 1;
  ram[819]  = 1;
  ram[820]  = 1;
  ram[821]  = 1;
  ram[822]  = 1;
  ram[823]  = 1;
  ram[824]  = 1;
  ram[825]  = 1;
  ram[826]  = 1;
  ram[827]  = 1;
  ram[828]  = 1;
  ram[829]  = 1;
  ram[830]  = 1;
  ram[831]  = 1;
  ram[832]  = 1;
  ram[833]  = 1;
  ram[834]  = 1;
  ram[835]  = 1;
  ram[836]  = 1;
  ram[837]  = 1;
  ram[838]  = 1;
  ram[839]  = 1;
  ram[840]  = 1;
  ram[841]  = 1;
  ram[842]  = 1;
  ram[843]  = 1;
  ram[844]  = 1;
  ram[845]  = 1;
  ram[846]  = 1;
  ram[847]  = 1;
  ram[848]  = 1;
  ram[849]  = 1;
  ram[850]  = 1;
  ram[851]  = 1;
  ram[852]  = 1;
  ram[853]  = 1;
  ram[854]  = 1;
  ram[855]  = 1;
  ram[856]  = 1;
  ram[857]  = 1;
  ram[858]  = 1;
  ram[859]  = 1;
  ram[860]  = 1;
  ram[861]  = 1;
  ram[862]  = 1;
  ram[863]  = 1;
  ram[864]  = 1;
  ram[865]  = 1;
  ram[866]  = 1;
  ram[867]  = 1;
  ram[868]  = 1;
  ram[869]  = 1;
  ram[870]  = 1;
  ram[871]  = 1;
  ram[872]  = 1;
  ram[873]  = 1;
  ram[874]  = 1;
  ram[875]  = 1;
  ram[876]  = 1;
  ram[877]  = 1;
  ram[878]  = 1;
  ram[879]  = 1;
  ram[880]  = 1;
  ram[881]  = 1;
  ram[882]  = 1;
  ram[883]  = 1;
  ram[884]  = 1;
  ram[885]  = 1;
  ram[886]  = 1;
  ram[887]  = 1;
  ram[888]  = 1;
  ram[889]  = 1;
  ram[890]  = 1;
  ram[891]  = 1;
  ram[892]  = 1;
  ram[893]  = 1;
  ram[894]  = 1;
  ram[895]  = 1;
  ram[896]  = 1;
  ram[897]  = 1;
  ram[898]  = 1;
  ram[899]  = 1;
  ram[900]  = 1;
  ram[901]  = 1;
  ram[902]  = 1;
  ram[903]  = 1;
  ram[904]  = 1;
  ram[905]  = 1;
  ram[906]  = 1;
  ram[907]  = 1;
  ram[908]  = 1;
  ram[909]  = 1;
  ram[910]  = 1;
  ram[911]  = 1;
  ram[912]  = 1;
  ram[913]  = 1;
  ram[914]  = 1;
  ram[915]  = 1;
  ram[916]  = 1;
  ram[917]  = 1;
  ram[918]  = 1;
  ram[919]  = 1;
  ram[920]  = 1;
  ram[921]  = 1;
  ram[922]  = 1;
  ram[923]  = 1;
  ram[924]  = 1;
  ram[925]  = 1;
  ram[926]  = 1;
  ram[927]  = 1;
  ram[928]  = 1;
  ram[929]  = 1;
  ram[930]  = 1;
  ram[931]  = 1;
  ram[932]  = 1;
  ram[933]  = 1;
  ram[934]  = 1;
  ram[935]  = 1;
  ram[936]  = 1;
  ram[937]  = 1;
  ram[938]  = 1;
  ram[939]  = 1;
  ram[940]  = 1;
  ram[941]  = 1;
  ram[942]  = 1;
  ram[943]  = 1;
  ram[944]  = 1;
  ram[945]  = 1;
  ram[946]  = 1;
  ram[947]  = 1;
  ram[948]  = 1;
  ram[949]  = 1;
  ram[950]  = 1;
  ram[951]  = 1;
  ram[952]  = 1;
  ram[953]  = 1;
  ram[954]  = 1;
  ram[955]  = 1;
  ram[956]  = 1;
  ram[957]  = 1;
  ram[958]  = 1;
  ram[959]  = 1;
  ram[960]  = 1;
  ram[961]  = 1;
  ram[962]  = 1;
  ram[963]  = 1;
  ram[964]  = 1;
  ram[965]  = 1;
  ram[966]  = 1;
  ram[967]  = 1;
  ram[968]  = 1;
  ram[969]  = 1;
  ram[970]  = 1;
  ram[971]  = 1;
  ram[972]  = 1;
  ram[973]  = 1;
  ram[974]  = 1;
  ram[975]  = 1;
  ram[976]  = 1;
  ram[977]  = 1;
  ram[978]  = 1;
  ram[979]  = 1;
  ram[980]  = 1;
  ram[981]  = 1;
  ram[982]  = 1;
  ram[983]  = 1;
  ram[984]  = 1;
  ram[985]  = 1;
  ram[986]  = 1;
  ram[987]  = 1;
  ram[988]  = 1;
  ram[989]  = 1;
  ram[990]  = 1;
  ram[991]  = 1;
  ram[992]  = 1;
  ram[993]  = 1;
  ram[994]  = 1;
  ram[995]  = 1;
  ram[996]  = 1;
  ram[997]  = 1;
  ram[998]  = 1;
  ram[999]  = 1;
  ram[1000]  = 1;
  ram[1001]  = 1;
  ram[1002]  = 1;
  ram[1003]  = 1;
  ram[1004]  = 1;
  ram[1005]  = 1;
  ram[1006]  = 1;
  ram[1007]  = 1;
  ram[1008]  = 1;
  ram[1009]  = 1;
  ram[1010]  = 1;
  ram[1011]  = 1;
  ram[1012]  = 1;
  ram[1013]  = 1;
  ram[1014]  = 1;
  ram[1015]  = 1;
  ram[1016]  = 1;
  ram[1017]  = 1;
  ram[1018]  = 1;
  ram[1019]  = 1;
  ram[1020]  = 1;
  ram[1021]  = 1;
  ram[1022]  = 1;
  ram[1023]  = 1;
  ram[1024]  = 1;
  ram[1025]  = 1;
  ram[1026]  = 1;
  ram[1027]  = 1;
  ram[1028]  = 1;
  ram[1029]  = 1;
  ram[1030]  = 1;
  ram[1031]  = 1;
  ram[1032]  = 1;
  ram[1033]  = 1;
  ram[1034]  = 1;
  ram[1035]  = 1;
  ram[1036]  = 1;
  ram[1037]  = 1;
  ram[1038]  = 1;
  ram[1039]  = 1;
  ram[1040]  = 1;
  ram[1041]  = 1;
  ram[1042]  = 1;
  ram[1043]  = 1;
  ram[1044]  = 1;
  ram[1045]  = 1;
  ram[1046]  = 1;
  ram[1047]  = 1;
  ram[1048]  = 1;
  ram[1049]  = 1;
  ram[1050]  = 1;
  ram[1051]  = 1;
  ram[1052]  = 1;
  ram[1053]  = 1;
  ram[1054]  = 1;
  ram[1055]  = 1;
  ram[1056]  = 1;
  ram[1057]  = 1;
  ram[1058]  = 1;
  ram[1059]  = 1;
  ram[1060]  = 1;
  ram[1061]  = 1;
  ram[1062]  = 1;
  ram[1063]  = 1;
  ram[1064]  = 1;
  ram[1065]  = 1;
  ram[1066]  = 1;
  ram[1067]  = 1;
  ram[1068]  = 1;
  ram[1069]  = 1;
  ram[1070]  = 1;
  ram[1071]  = 1;
  ram[1072]  = 1;
  ram[1073]  = 1;
  ram[1074]  = 1;
  ram[1075]  = 1;
  ram[1076]  = 1;
  ram[1077]  = 1;
  ram[1078]  = 1;
  ram[1079]  = 1;
  ram[1080]  = 1;
  ram[1081]  = 1;
  ram[1082]  = 1;
  ram[1083]  = 1;
  ram[1084]  = 1;
  ram[1085]  = 1;
  ram[1086]  = 1;
  ram[1087]  = 1;
  ram[1088]  = 1;
  ram[1089]  = 1;
  ram[1090]  = 1;
  ram[1091]  = 1;
  ram[1092]  = 1;
  ram[1093]  = 1;
  ram[1094]  = 1;
  ram[1095]  = 1;
  ram[1096]  = 1;
  ram[1097]  = 1;
  ram[1098]  = 1;
  ram[1099]  = 1;
  ram[1100]  = 1;
  ram[1101]  = 1;
  ram[1102]  = 1;
  ram[1103]  = 1;
  ram[1104]  = 1;
  ram[1105]  = 1;
  ram[1106]  = 1;
  ram[1107]  = 1;
  ram[1108]  = 1;
  ram[1109]  = 1;
  ram[1110]  = 1;
  ram[1111]  = 1;
  ram[1112]  = 1;
  ram[1113]  = 1;
  ram[1114]  = 1;
  ram[1115]  = 1;
  ram[1116]  = 1;
  ram[1117]  = 1;
  ram[1118]  = 1;
  ram[1119]  = 1;
  ram[1120]  = 1;
  ram[1121]  = 1;
  ram[1122]  = 1;
  ram[1123]  = 1;
  ram[1124]  = 1;
  ram[1125]  = 1;
  ram[1126]  = 1;
  ram[1127]  = 1;
  ram[1128]  = 1;
  ram[1129]  = 1;
  ram[1130]  = 1;
  ram[1131]  = 1;
  ram[1132]  = 1;
  ram[1133]  = 1;
  ram[1134]  = 1;
  ram[1135]  = 1;
  ram[1136]  = 1;
  ram[1137]  = 1;
  ram[1138]  = 1;
  ram[1139]  = 1;
  ram[1140]  = 1;
  ram[1141]  = 1;
  ram[1142]  = 1;
  ram[1143]  = 1;
  ram[1144]  = 1;
  ram[1145]  = 1;
  ram[1146]  = 1;
  ram[1147]  = 1;
  ram[1148]  = 1;
  ram[1149]  = 1;
  ram[1150]  = 1;
  ram[1151]  = 1;
  ram[1152]  = 1;
  ram[1153]  = 1;
  ram[1154]  = 1;
  ram[1155]  = 1;
  ram[1156]  = 1;
  ram[1157]  = 1;
  ram[1158]  = 1;
  ram[1159]  = 1;
  ram[1160]  = 1;
  ram[1161]  = 1;
  ram[1162]  = 1;
  ram[1163]  = 1;
  ram[1164]  = 1;
  ram[1165]  = 1;
  ram[1166]  = 1;
  ram[1167]  = 1;
  ram[1168]  = 1;
  ram[1169]  = 1;
  ram[1170]  = 1;
  ram[1171]  = 1;
  ram[1172]  = 1;
  ram[1173]  = 1;
  ram[1174]  = 1;
  ram[1175]  = 1;
  ram[1176]  = 1;
  ram[1177]  = 1;
  ram[1178]  = 1;
  ram[1179]  = 1;
  ram[1180]  = 1;
  ram[1181]  = 1;
  ram[1182]  = 1;
  ram[1183]  = 1;
  ram[1184]  = 1;
  ram[1185]  = 1;
  ram[1186]  = 1;
  ram[1187]  = 1;
  ram[1188]  = 1;
  ram[1189]  = 1;
  ram[1190]  = 1;
  ram[1191]  = 1;
  ram[1192]  = 1;
  ram[1193]  = 1;
  ram[1194]  = 1;
  ram[1195]  = 1;
  ram[1196]  = 1;
  ram[1197]  = 1;
  ram[1198]  = 1;
  ram[1199]  = 1;
  ram[1200]  = 1;
  ram[1201]  = 1;
  ram[1202]  = 1;
  ram[1203]  = 1;
  ram[1204]  = 1;
  ram[1205]  = 1;
  ram[1206]  = 1;
  ram[1207]  = 1;
  ram[1208]  = 1;
  ram[1209]  = 1;
  ram[1210]  = 1;
  ram[1211]  = 1;
  ram[1212]  = 1;
  ram[1213]  = 1;
  ram[1214]  = 1;
  ram[1215]  = 1;
  ram[1216]  = 1;
  ram[1217]  = 1;
  ram[1218]  = 1;
  ram[1219]  = 1;
  ram[1220]  = 1;
  ram[1221]  = 1;
  ram[1222]  = 1;
  ram[1223]  = 1;
  ram[1224]  = 1;
  ram[1225]  = 1;
  ram[1226]  = 1;
  ram[1227]  = 1;
  ram[1228]  = 1;
  ram[1229]  = 1;
  ram[1230]  = 1;
  ram[1231]  = 1;
  ram[1232]  = 1;
  ram[1233]  = 1;
  ram[1234]  = 1;
  ram[1235]  = 1;
  ram[1236]  = 1;
  ram[1237]  = 1;
  ram[1238]  = 1;
  ram[1239]  = 1;
  ram[1240]  = 1;
  ram[1241]  = 1;
  ram[1242]  = 1;
  ram[1243]  = 1;
  ram[1244]  = 1;
  ram[1245]  = 1;
  ram[1246]  = 1;
  ram[1247]  = 1;
  ram[1248]  = 1;
  ram[1249]  = 1;
  ram[1250]  = 1;
  ram[1251]  = 1;
  ram[1252]  = 1;
  ram[1253]  = 1;
  ram[1254]  = 1;
  ram[1255]  = 1;
  ram[1256]  = 1;
  ram[1257]  = 1;
  ram[1258]  = 1;
  ram[1259]  = 1;
  ram[1260]  = 1;
  ram[1261]  = 1;
  ram[1262]  = 1;
  ram[1263]  = 1;
  ram[1264]  = 1;
  ram[1265]  = 1;
  ram[1266]  = 1;
  ram[1267]  = 1;
  ram[1268]  = 1;
  ram[1269]  = 1;
  ram[1270]  = 1;
  ram[1271]  = 1;
  ram[1272]  = 1;
  ram[1273]  = 1;
  ram[1274]  = 1;
  ram[1275]  = 1;
  ram[1276]  = 1;
  ram[1277]  = 1;
  ram[1278]  = 1;
  ram[1279]  = 1;
  ram[1280]  = 1;
  ram[1281]  = 1;
  ram[1282]  = 1;
  ram[1283]  = 1;
  ram[1284]  = 1;
  ram[1285]  = 1;
  ram[1286]  = 1;
  ram[1287]  = 1;
  ram[1288]  = 1;
  ram[1289]  = 1;
  ram[1290]  = 1;
  ram[1291]  = 1;
  ram[1292]  = 1;
  ram[1293]  = 1;
  ram[1294]  = 1;
  ram[1295]  = 1;
  ram[1296]  = 1;
  ram[1297]  = 1;
  ram[1298]  = 1;
  ram[1299]  = 1;
  ram[1300]  = 1;
  ram[1301]  = 1;
  ram[1302]  = 1;
  ram[1303]  = 1;
  ram[1304]  = 1;
  ram[1305]  = 1;
  ram[1306]  = 1;
  ram[1307]  = 1;
  ram[1308]  = 1;
  ram[1309]  = 1;
  ram[1310]  = 1;
  ram[1311]  = 1;
  ram[1312]  = 1;
  ram[1313]  = 1;
  ram[1314]  = 1;
  ram[1315]  = 1;
  ram[1316]  = 1;
  ram[1317]  = 1;
  ram[1318]  = 1;
  ram[1319]  = 1;
  ram[1320]  = 1;
  ram[1321]  = 1;
  ram[1322]  = 1;
  ram[1323]  = 1;
  ram[1324]  = 1;
  ram[1325]  = 1;
  ram[1326]  = 1;
  ram[1327]  = 1;
  ram[1328]  = 1;
  ram[1329]  = 1;
  ram[1330]  = 1;
  ram[1331]  = 1;
  ram[1332]  = 1;
  ram[1333]  = 1;
  ram[1334]  = 1;
  ram[1335]  = 1;
  ram[1336]  = 1;
  ram[1337]  = 1;
  ram[1338]  = 1;
  ram[1339]  = 1;
  ram[1340]  = 1;
  ram[1341]  = 1;
  ram[1342]  = 1;
  ram[1343]  = 1;
  ram[1344]  = 1;
  ram[1345]  = 1;
  ram[1346]  = 1;
  ram[1347]  = 1;
  ram[1348]  = 1;
  ram[1349]  = 1;
  ram[1350]  = 1;
  ram[1351]  = 1;
  ram[1352]  = 1;
  ram[1353]  = 1;
  ram[1354]  = 1;
  ram[1355]  = 1;
  ram[1356]  = 1;
  ram[1357]  = 1;
  ram[1358]  = 1;
  ram[1359]  = 1;
  ram[1360]  = 1;
  ram[1361]  = 1;
  ram[1362]  = 1;
  ram[1363]  = 1;
  ram[1364]  = 1;
  ram[1365]  = 1;
  ram[1366]  = 1;
  ram[1367]  = 1;
  ram[1368]  = 1;
  ram[1369]  = 1;
  ram[1370]  = 1;
  ram[1371]  = 1;
  ram[1372]  = 1;
  ram[1373]  = 1;
  ram[1374]  = 1;
  ram[1375]  = 1;
  ram[1376]  = 1;
  ram[1377]  = 1;
  ram[1378]  = 1;
  ram[1379]  = 1;
  ram[1380]  = 1;
  ram[1381]  = 1;
  ram[1382]  = 1;
  ram[1383]  = 1;
  ram[1384]  = 1;
  ram[1385]  = 1;
  ram[1386]  = 1;
  ram[1387]  = 1;
  ram[1388]  = 1;
  ram[1389]  = 1;
  ram[1390]  = 1;
  ram[1391]  = 1;
  ram[1392]  = 1;
  ram[1393]  = 1;
  ram[1394]  = 1;
  ram[1395]  = 1;
  ram[1396]  = 1;
  ram[1397]  = 1;
  ram[1398]  = 1;
  ram[1399]  = 1;
  ram[1400]  = 1;
  ram[1401]  = 1;
  ram[1402]  = 1;
  ram[1403]  = 1;
  ram[1404]  = 1;
  ram[1405]  = 1;
  ram[1406]  = 1;
  ram[1407]  = 1;
  ram[1408]  = 1;
  ram[1409]  = 1;
  ram[1410]  = 1;
  ram[1411]  = 1;
  ram[1412]  = 1;
  ram[1413]  = 1;
  ram[1414]  = 1;
  ram[1415]  = 1;
  ram[1416]  = 1;
  ram[1417]  = 1;
  ram[1418]  = 1;
  ram[1419]  = 1;
  ram[1420]  = 1;
  ram[1421]  = 1;
  ram[1422]  = 1;
  ram[1423]  = 1;
  ram[1424]  = 1;
  ram[1425]  = 1;
  ram[1426]  = 1;
  ram[1427]  = 1;
  ram[1428]  = 1;
  ram[1429]  = 1;
  ram[1430]  = 1;
  ram[1431]  = 1;
  ram[1432]  = 1;
  ram[1433]  = 1;
  ram[1434]  = 1;
  ram[1435]  = 1;
  ram[1436]  = 1;
  ram[1437]  = 1;
  ram[1438]  = 1;
  ram[1439]  = 1;
  ram[1440]  = 1;
  ram[1441]  = 1;
  ram[1442]  = 1;
  ram[1443]  = 1;
  ram[1444]  = 1;
  ram[1445]  = 1;
  ram[1446]  = 1;
  ram[1447]  = 1;
  ram[1448]  = 1;
  ram[1449]  = 1;
  ram[1450]  = 1;
  ram[1451]  = 1;
  ram[1452]  = 1;
  ram[1453]  = 1;
  ram[1454]  = 1;
  ram[1455]  = 1;
  ram[1456]  = 1;
  ram[1457]  = 1;
  ram[1458]  = 1;
  ram[1459]  = 1;
  ram[1460]  = 1;
  ram[1461]  = 1;
  ram[1462]  = 1;
  ram[1463]  = 1;
  ram[1464]  = 1;
  ram[1465]  = 1;
  ram[1466]  = 1;
  ram[1467]  = 1;
  ram[1468]  = 1;
  ram[1469]  = 1;
  ram[1470]  = 1;
  ram[1471]  = 1;
  ram[1472]  = 1;
  ram[1473]  = 1;
  ram[1474]  = 1;
  ram[1475]  = 1;
  ram[1476]  = 1;
  ram[1477]  = 1;
  ram[1478]  = 1;
  ram[1479]  = 1;
  ram[1480]  = 1;
  ram[1481]  = 1;
  ram[1482]  = 1;
  ram[1483]  = 1;
  ram[1484]  = 1;
  ram[1485]  = 1;
  ram[1486]  = 1;
  ram[1487]  = 1;
  ram[1488]  = 1;
  ram[1489]  = 1;
  ram[1490]  = 1;
  ram[1491]  = 1;
  ram[1492]  = 1;
  ram[1493]  = 1;
  ram[1494]  = 1;
  ram[1495]  = 1;
  ram[1496]  = 1;
  ram[1497]  = 1;
  ram[1498]  = 1;
  ram[1499]  = 1;
  ram[1500]  = 1;
  ram[1501]  = 1;
  ram[1502]  = 1;
  ram[1503]  = 1;
  ram[1504]  = 1;
  ram[1505]  = 1;
  ram[1506]  = 1;
  ram[1507]  = 1;
  ram[1508]  = 1;
  ram[1509]  = 1;
  ram[1510]  = 1;
  ram[1511]  = 1;
  ram[1512]  = 1;
  ram[1513]  = 1;
  ram[1514]  = 1;
  ram[1515]  = 1;
  ram[1516]  = 1;
  ram[1517]  = 1;
  ram[1518]  = 1;
  ram[1519]  = 1;
  ram[1520]  = 1;
  ram[1521]  = 1;
  ram[1522]  = 1;
  ram[1523]  = 1;
  ram[1524]  = 1;
  ram[1525]  = 1;
  ram[1526]  = 1;
  ram[1527]  = 1;
  ram[1528]  = 1;
  ram[1529]  = 1;
  ram[1530]  = 1;
  ram[1531]  = 1;
  ram[1532]  = 1;
  ram[1533]  = 1;
  ram[1534]  = 1;
  ram[1535]  = 1;
  ram[1536]  = 1;
  ram[1537]  = 1;
  ram[1538]  = 1;
  ram[1539]  = 1;
  ram[1540]  = 1;
  ram[1541]  = 1;
  ram[1542]  = 1;
  ram[1543]  = 1;
  ram[1544]  = 1;
  ram[1545]  = 1;
  ram[1546]  = 1;
  ram[1547]  = 1;
  ram[1548]  = 1;
  ram[1549]  = 1;
  ram[1550]  = 1;
  ram[1551]  = 1;
  ram[1552]  = 1;
  ram[1553]  = 1;
  ram[1554]  = 1;
  ram[1555]  = 1;
  ram[1556]  = 1;
  ram[1557]  = 1;
  ram[1558]  = 1;
  ram[1559]  = 1;
  ram[1560]  = 1;
  ram[1561]  = 1;
  ram[1562]  = 1;
  ram[1563]  = 1;
  ram[1564]  = 1;
  ram[1565]  = 1;
  ram[1566]  = 1;
  ram[1567]  = 1;
  ram[1568]  = 1;
  ram[1569]  = 1;
  ram[1570]  = 1;
  ram[1571]  = 1;
  ram[1572]  = 1;
  ram[1573]  = 1;
  ram[1574]  = 1;
  ram[1575]  = 1;
  ram[1576]  = 1;
  ram[1577]  = 1;
  ram[1578]  = 1;
  ram[1579]  = 1;
  ram[1580]  = 1;
  ram[1581]  = 1;
  ram[1582]  = 1;
  ram[1583]  = 1;
  ram[1584]  = 1;
  ram[1585]  = 1;
  ram[1586]  = 1;
  ram[1587]  = 1;
  ram[1588]  = 1;
  ram[1589]  = 1;
  ram[1590]  = 1;
  ram[1591]  = 1;
  ram[1592]  = 1;
  ram[1593]  = 1;
  ram[1594]  = 1;
  ram[1595]  = 1;
  ram[1596]  = 1;
  ram[1597]  = 1;
  ram[1598]  = 1;
  ram[1599]  = 1;
  ram[1600]  = 1;
  ram[1601]  = 1;
  ram[1602]  = 1;
  ram[1603]  = 1;
  ram[1604]  = 1;
  ram[1605]  = 1;
  ram[1606]  = 1;
  ram[1607]  = 1;
  ram[1608]  = 1;
  ram[1609]  = 1;
  ram[1610]  = 1;
  ram[1611]  = 1;
  ram[1612]  = 1;
  ram[1613]  = 1;
  ram[1614]  = 1;
  ram[1615]  = 1;
  ram[1616]  = 1;
  ram[1617]  = 1;
  ram[1618]  = 1;
  ram[1619]  = 1;
  ram[1620]  = 1;
  ram[1621]  = 1;
  ram[1622]  = 1;
  ram[1623]  = 1;
  ram[1624]  = 1;
  ram[1625]  = 1;
  ram[1626]  = 1;
  ram[1627]  = 1;
  ram[1628]  = 1;
  ram[1629]  = 1;
  ram[1630]  = 1;
  ram[1631]  = 1;
  ram[1632]  = 1;
  ram[1633]  = 1;
  ram[1634]  = 1;
  ram[1635]  = 1;
  ram[1636]  = 1;
  ram[1637]  = 1;
  ram[1638]  = 1;
  ram[1639]  = 1;
  ram[1640]  = 1;
  ram[1641]  = 1;
  ram[1642]  = 1;
  ram[1643]  = 1;
  ram[1644]  = 1;
  ram[1645]  = 1;
  ram[1646]  = 1;
  ram[1647]  = 1;
  ram[1648]  = 1;
  ram[1649]  = 1;
  ram[1650]  = 1;
  ram[1651]  = 1;
  ram[1652]  = 1;
  ram[1653]  = 1;
  ram[1654]  = 1;
  ram[1655]  = 1;
  ram[1656]  = 1;
  ram[1657]  = 1;
  ram[1658]  = 1;
  ram[1659]  = 1;
  ram[1660]  = 1;
  ram[1661]  = 1;
  ram[1662]  = 1;
  ram[1663]  = 1;
  ram[1664]  = 1;
  ram[1665]  = 1;
  ram[1666]  = 1;
  ram[1667]  = 1;
  ram[1668]  = 1;
  ram[1669]  = 1;
  ram[1670]  = 1;
  ram[1671]  = 1;
  ram[1672]  = 1;
  ram[1673]  = 1;
  ram[1674]  = 1;
  ram[1675]  = 1;
  ram[1676]  = 1;
  ram[1677]  = 1;
  ram[1678]  = 1;
  ram[1679]  = 1;
  ram[1680]  = 1;
  ram[1681]  = 1;
  ram[1682]  = 1;
  ram[1683]  = 1;
  ram[1684]  = 1;
  ram[1685]  = 1;
  ram[1686]  = 1;
  ram[1687]  = 1;
  ram[1688]  = 1;
  ram[1689]  = 1;
  ram[1690]  = 1;
  ram[1691]  = 1;
  ram[1692]  = 1;
  ram[1693]  = 1;
  ram[1694]  = 1;
  ram[1695]  = 1;
  ram[1696]  = 1;
  ram[1697]  = 1;
  ram[1698]  = 1;
  ram[1699]  = 1;
  ram[1700]  = 1;
  ram[1701]  = 1;
  ram[1702]  = 1;
  ram[1703]  = 1;
  ram[1704]  = 1;
  ram[1705]  = 1;
  ram[1706]  = 1;
  ram[1707]  = 1;
  ram[1708]  = 1;
  ram[1709]  = 1;
  ram[1710]  = 1;
  ram[1711]  = 1;
  ram[1712]  = 1;
  ram[1713]  = 1;
  ram[1714]  = 1;
  ram[1715]  = 1;
  ram[1716]  = 1;
  ram[1717]  = 1;
  ram[1718]  = 1;
  ram[1719]  = 1;
  ram[1720]  = 1;
  ram[1721]  = 1;
  ram[1722]  = 1;
  ram[1723]  = 1;
  ram[1724]  = 1;
  ram[1725]  = 1;
  ram[1726]  = 1;
  ram[1727]  = 1;
  ram[1728]  = 1;
  ram[1729]  = 1;
  ram[1730]  = 1;
  ram[1731]  = 1;
  ram[1732]  = 1;
  ram[1733]  = 1;
  ram[1734]  = 1;
  ram[1735]  = 1;
  ram[1736]  = 1;
  ram[1737]  = 1;
  ram[1738]  = 1;
  ram[1739]  = 1;
  ram[1740]  = 1;
  ram[1741]  = 1;
  ram[1742]  = 1;
  ram[1743]  = 1;
  ram[1744]  = 1;
  ram[1745]  = 1;
  ram[1746]  = 1;
  ram[1747]  = 1;
  ram[1748]  = 1;
  ram[1749]  = 1;
  ram[1750]  = 1;
  ram[1751]  = 1;
  ram[1752]  = 1;
  ram[1753]  = 1;
  ram[1754]  = 1;
  ram[1755]  = 1;
  ram[1756]  = 1;
  ram[1757]  = 1;
  ram[1758]  = 1;
  ram[1759]  = 1;
  ram[1760]  = 1;
  ram[1761]  = 1;
  ram[1762]  = 1;
  ram[1763]  = 1;
  ram[1764]  = 1;
  ram[1765]  = 1;
  ram[1766]  = 1;
  ram[1767]  = 1;
  ram[1768]  = 1;
  ram[1769]  = 1;
  ram[1770]  = 1;
  ram[1771]  = 1;
  ram[1772]  = 1;
  ram[1773]  = 1;
  ram[1774]  = 1;
  ram[1775]  = 1;
  ram[1776]  = 1;
  ram[1777]  = 1;
  ram[1778]  = 1;
  ram[1779]  = 1;
  ram[1780]  = 1;
  ram[1781]  = 1;
  ram[1782]  = 1;
  ram[1783]  = 1;
  ram[1784]  = 1;
  ram[1785]  = 1;
  ram[1786]  = 1;
  ram[1787]  = 1;
  ram[1788]  = 1;
  ram[1789]  = 1;
  ram[1790]  = 1;
  ram[1791]  = 1;
  ram[1792]  = 1;
  ram[1793]  = 1;
  ram[1794]  = 1;
  ram[1795]  = 1;
  ram[1796]  = 1;
  ram[1797]  = 1;
  ram[1798]  = 1;
  ram[1799]  = 1;
  ram[1800]  = 1;
  ram[1801]  = 1;
  ram[1802]  = 1;
  ram[1803]  = 1;
  ram[1804]  = 1;
  ram[1805]  = 1;
  ram[1806]  = 1;
  ram[1807]  = 1;
  ram[1808]  = 1;
  ram[1809]  = 1;
  ram[1810]  = 1;
  ram[1811]  = 1;
  ram[1812]  = 1;
  ram[1813]  = 1;
  ram[1814]  = 1;
  ram[1815]  = 1;
  ram[1816]  = 1;
  ram[1817]  = 1;
  ram[1818]  = 1;
  ram[1819]  = 1;
  ram[1820]  = 1;
  ram[1821]  = 1;
  ram[1822]  = 1;
  ram[1823]  = 1;
  ram[1824]  = 1;
  ram[1825]  = 1;
  ram[1826]  = 1;
  ram[1827]  = 1;
  ram[1828]  = 1;
  ram[1829]  = 1;
  ram[1830]  = 1;
  ram[1831]  = 1;
  ram[1832]  = 1;
  ram[1833]  = 1;
  ram[1834]  = 1;
  ram[1835]  = 1;
  ram[1836]  = 1;
  ram[1837]  = 1;
  ram[1838]  = 1;
  ram[1839]  = 1;
  ram[1840]  = 1;
  ram[1841]  = 1;
  ram[1842]  = 1;
  ram[1843]  = 1;
  ram[1844]  = 1;
  ram[1845]  = 1;
  ram[1846]  = 1;
  ram[1847]  = 1;
  ram[1848]  = 1;
  ram[1849]  = 1;
  ram[1850]  = 1;
  ram[1851]  = 1;
  ram[1852]  = 1;
  ram[1853]  = 1;
  ram[1854]  = 1;
  ram[1855]  = 1;
  ram[1856]  = 1;
  ram[1857]  = 1;
  ram[1858]  = 1;
  ram[1859]  = 1;
  ram[1860]  = 1;
  ram[1861]  = 1;
  ram[1862]  = 1;
  ram[1863]  = 1;
  ram[1864]  = 1;
  ram[1865]  = 1;
  ram[1866]  = 1;
  ram[1867]  = 1;
  ram[1868]  = 1;
  ram[1869]  = 1;
  ram[1870]  = 1;
  ram[1871]  = 1;
  ram[1872]  = 1;
  ram[1873]  = 1;
  ram[1874]  = 1;
  ram[1875]  = 1;
  ram[1876]  = 1;
  ram[1877]  = 1;
  ram[1878]  = 1;
  ram[1879]  = 1;
  ram[1880]  = 1;
  ram[1881]  = 1;
  ram[1882]  = 1;
  ram[1883]  = 1;
  ram[1884]  = 1;
  ram[1885]  = 1;
  ram[1886]  = 1;
  ram[1887]  = 1;
  ram[1888]  = 1;
  ram[1889]  = 1;
  ram[1890]  = 1;
  ram[1891]  = 1;
  ram[1892]  = 1;
  ram[1893]  = 1;
  ram[1894]  = 1;
  ram[1895]  = 1;
  ram[1896]  = 1;
  ram[1897]  = 1;
  ram[1898]  = 1;
  ram[1899]  = 1;
  ram[1900]  = 1;
  ram[1901]  = 1;
  ram[1902]  = 1;
  ram[1903]  = 1;
  ram[1904]  = 1;
  ram[1905]  = 1;
  ram[1906]  = 1;
  ram[1907]  = 1;
  ram[1908]  = 1;
  ram[1909]  = 1;
  ram[1910]  = 1;
  ram[1911]  = 1;
  ram[1912]  = 1;
  ram[1913]  = 1;
  ram[1914]  = 1;
  ram[1915]  = 1;
  ram[1916]  = 1;
  ram[1917]  = 1;
  ram[1918]  = 1;
  ram[1919]  = 1;
  ram[1920]  = 1;
  ram[1921]  = 1;
  ram[1922]  = 1;
  ram[1923]  = 1;
  ram[1924]  = 1;
  ram[1925]  = 1;
  ram[1926]  = 1;
  ram[1927]  = 1;
  ram[1928]  = 1;
  ram[1929]  = 1;
  ram[1930]  = 1;
  ram[1931]  = 1;
  ram[1932]  = 1;
  ram[1933]  = 1;
  ram[1934]  = 1;
  ram[1935]  = 1;
  ram[1936]  = 1;
  ram[1937]  = 1;
  ram[1938]  = 1;
  ram[1939]  = 1;
  ram[1940]  = 1;
  ram[1941]  = 1;
  ram[1942]  = 1;
  ram[1943]  = 1;
  ram[1944]  = 1;
  ram[1945]  = 1;
  ram[1946]  = 1;
  ram[1947]  = 1;
  ram[1948]  = 1;
  ram[1949]  = 1;
  ram[1950]  = 1;
  ram[1951]  = 1;
  ram[1952]  = 1;
  ram[1953]  = 1;
  ram[1954]  = 1;
  ram[1955]  = 1;
  ram[1956]  = 1;
  ram[1957]  = 1;
  ram[1958]  = 1;
  ram[1959]  = 1;
  ram[1960]  = 1;
  ram[1961]  = 1;
  ram[1962]  = 1;
  ram[1963]  = 1;
  ram[1964]  = 1;
  ram[1965]  = 1;
  ram[1966]  = 1;
  ram[1967]  = 1;
  ram[1968]  = 1;
  ram[1969]  = 1;
  ram[1970]  = 1;
  ram[1971]  = 1;
  ram[1972]  = 1;
  ram[1973]  = 1;
  ram[1974]  = 1;
  ram[1975]  = 1;
  ram[1976]  = 1;
  ram[1977]  = 1;
  ram[1978]  = 1;
  ram[1979]  = 1;
  ram[1980]  = 1;
  ram[1981]  = 1;
  ram[1982]  = 1;
  ram[1983]  = 1;
  ram[1984]  = 1;
  ram[1985]  = 1;
  ram[1986]  = 1;
  ram[1987]  = 1;
  ram[1988]  = 1;
  ram[1989]  = 1;
  ram[1990]  = 1;
  ram[1991]  = 1;
  ram[1992]  = 1;
  ram[1993]  = 1;
  ram[1994]  = 1;
  ram[1995]  = 1;
  ram[1996]  = 1;
  ram[1997]  = 1;
  ram[1998]  = 1;
  ram[1999]  = 1;
  ram[2000]  = 1;
  ram[2001]  = 1;
  ram[2002]  = 1;
  ram[2003]  = 1;
  ram[2004]  = 1;
  ram[2005]  = 1;
  ram[2006]  = 1;
  ram[2007]  = 1;
  ram[2008]  = 1;
  ram[2009]  = 1;
  ram[2010]  = 1;
  ram[2011]  = 1;
  ram[2012]  = 1;
  ram[2013]  = 1;
  ram[2014]  = 1;
  ram[2015]  = 1;
  ram[2016]  = 1;
  ram[2017]  = 1;
  ram[2018]  = 1;
  ram[2019]  = 1;
  ram[2020]  = 1;
  ram[2021]  = 1;
  ram[2022]  = 1;
  ram[2023]  = 1;
  ram[2024]  = 1;
  ram[2025]  = 1;
  ram[2026]  = 1;
  ram[2027]  = 1;
  ram[2028]  = 1;
  ram[2029]  = 1;
  ram[2030]  = 1;
  ram[2031]  = 1;
  ram[2032]  = 1;
  ram[2033]  = 1;
  ram[2034]  = 1;
  ram[2035]  = 1;
  ram[2036]  = 1;
  ram[2037]  = 1;
  ram[2038]  = 1;
  ram[2039]  = 1;
  ram[2040]  = 1;
  ram[2041]  = 1;
  ram[2042]  = 1;
  ram[2043]  = 1;
  ram[2044]  = 1;
  ram[2045]  = 1;
  ram[2046]  = 1;
  ram[2047]  = 1;
  ram[2048]  = 1;
  ram[2049]  = 1;
  ram[2050]  = 1;
  ram[2051]  = 1;
  ram[2052]  = 1;
  ram[2053]  = 1;
  ram[2054]  = 1;
  ram[2055]  = 1;
  ram[2056]  = 1;
  ram[2057]  = 1;
  ram[2058]  = 1;
  ram[2059]  = 1;
  ram[2060]  = 1;
  ram[2061]  = 1;
  ram[2062]  = 1;
  ram[2063]  = 1;
  ram[2064]  = 1;
  ram[2065]  = 1;
  ram[2066]  = 1;
  ram[2067]  = 1;
  ram[2068]  = 1;
  ram[2069]  = 1;
  ram[2070]  = 1;
  ram[2071]  = 1;
  ram[2072]  = 1;
  ram[2073]  = 1;
  ram[2074]  = 1;
  ram[2075]  = 1;
  ram[2076]  = 1;
  ram[2077]  = 1;
  ram[2078]  = 1;
  ram[2079]  = 1;
  ram[2080]  = 1;
  ram[2081]  = 1;
  ram[2082]  = 1;
  ram[2083]  = 1;
  ram[2084]  = 1;
  ram[2085]  = 1;
  ram[2086]  = 1;
  ram[2087]  = 1;
  ram[2088]  = 1;
  ram[2089]  = 1;
  ram[2090]  = 1;
  ram[2091]  = 1;
  ram[2092]  = 1;
  ram[2093]  = 1;
  ram[2094]  = 1;
  ram[2095]  = 1;
  ram[2096]  = 1;
  ram[2097]  = 1;
  ram[2098]  = 1;
  ram[2099]  = 1;
  ram[2100]  = 1;
  ram[2101]  = 1;
  ram[2102]  = 1;
  ram[2103]  = 1;
  ram[2104]  = 1;
  ram[2105]  = 1;
  ram[2106]  = 1;
  ram[2107]  = 1;
  ram[2108]  = 1;
  ram[2109]  = 1;
  ram[2110]  = 1;
  ram[2111]  = 1;
  ram[2112]  = 1;
  ram[2113]  = 1;
  ram[2114]  = 1;
  ram[2115]  = 1;
  ram[2116]  = 1;
  ram[2117]  = 1;
  ram[2118]  = 1;
  ram[2119]  = 1;
  ram[2120]  = 1;
  ram[2121]  = 1;
  ram[2122]  = 1;
  ram[2123]  = 1;
  ram[2124]  = 1;
  ram[2125]  = 1;
  ram[2126]  = 1;
  ram[2127]  = 1;
  ram[2128]  = 1;
  ram[2129]  = 1;
  ram[2130]  = 1;
  ram[2131]  = 1;
  ram[2132]  = 1;
  ram[2133]  = 1;
  ram[2134]  = 1;
  ram[2135]  = 1;
  ram[2136]  = 1;
  ram[2137]  = 1;
  ram[2138]  = 1;
  ram[2139]  = 1;
  ram[2140]  = 1;
  ram[2141]  = 1;
  ram[2142]  = 1;
  ram[2143]  = 1;
  ram[2144]  = 1;
  ram[2145]  = 1;
  ram[2146]  = 1;
  ram[2147]  = 1;
  ram[2148]  = 1;
  ram[2149]  = 1;
  ram[2150]  = 1;
  ram[2151]  = 1;
  ram[2152]  = 1;
  ram[2153]  = 1;
  ram[2154]  = 1;
  ram[2155]  = 1;
  ram[2156]  = 1;
  ram[2157]  = 1;
  ram[2158]  = 1;
  ram[2159]  = 1;
  ram[2160]  = 1;
  ram[2161]  = 1;
  ram[2162]  = 1;
  ram[2163]  = 1;
  ram[2164]  = 1;
  ram[2165]  = 1;
  ram[2166]  = 1;
  ram[2167]  = 1;
  ram[2168]  = 1;
  ram[2169]  = 1;
  ram[2170]  = 1;
  ram[2171]  = 1;
  ram[2172]  = 1;
  ram[2173]  = 1;
  ram[2174]  = 1;
  ram[2175]  = 1;
  ram[2176]  = 1;
  ram[2177]  = 1;
  ram[2178]  = 1;
  ram[2179]  = 1;
  ram[2180]  = 1;
  ram[2181]  = 1;
  ram[2182]  = 1;
  ram[2183]  = 1;
  ram[2184]  = 1;
  ram[2185]  = 1;
  ram[2186]  = 1;
  ram[2187]  = 1;
  ram[2188]  = 1;
  ram[2189]  = 1;
  ram[2190]  = 1;
  ram[2191]  = 1;
  ram[2192]  = 1;
  ram[2193]  = 1;
  ram[2194]  = 1;
  ram[2195]  = 1;
  ram[2196]  = 1;
  ram[2197]  = 1;
  ram[2198]  = 1;
  ram[2199]  = 1;
  ram[2200]  = 1;
  ram[2201]  = 1;
  ram[2202]  = 1;
  ram[2203]  = 1;
  ram[2204]  = 1;
  ram[2205]  = 1;
  ram[2206]  = 1;
  ram[2207]  = 1;
  ram[2208]  = 1;
  ram[2209]  = 1;
  ram[2210]  = 1;
  ram[2211]  = 1;
  ram[2212]  = 1;
  ram[2213]  = 1;
  ram[2214]  = 1;
  ram[2215]  = 1;
  ram[2216]  = 1;
  ram[2217]  = 1;
  ram[2218]  = 1;
  ram[2219]  = 1;
  ram[2220]  = 1;
  ram[2221]  = 1;
  ram[2222]  = 1;
  ram[2223]  = 1;
  ram[2224]  = 1;
  ram[2225]  = 1;
  ram[2226]  = 1;
  ram[2227]  = 1;
  ram[2228]  = 1;
  ram[2229]  = 1;
  ram[2230]  = 1;
  ram[2231]  = 1;
  ram[2232]  = 1;
  ram[2233]  = 1;
  ram[2234]  = 1;
  ram[2235]  = 1;
  ram[2236]  = 1;
  ram[2237]  = 1;
  ram[2238]  = 1;
  ram[2239]  = 1;
  ram[2240]  = 1;
  ram[2241]  = 1;
  ram[2242]  = 1;
  ram[2243]  = 1;
  ram[2244]  = 1;
  ram[2245]  = 1;
  ram[2246]  = 1;
  ram[2247]  = 1;
  ram[2248]  = 1;
  ram[2249]  = 1;
  ram[2250]  = 1;
  ram[2251]  = 1;
  ram[2252]  = 1;
  ram[2253]  = 1;
  ram[2254]  = 1;
  ram[2255]  = 1;
  ram[2256]  = 1;
  ram[2257]  = 1;
  ram[2258]  = 1;
  ram[2259]  = 1;
  ram[2260]  = 1;
  ram[2261]  = 1;
  ram[2262]  = 1;
  ram[2263]  = 1;
  ram[2264]  = 1;
  ram[2265]  = 1;
  ram[2266]  = 1;
  ram[2267]  = 1;
  ram[2268]  = 1;
  ram[2269]  = 1;
  ram[2270]  = 1;
  ram[2271]  = 1;
  ram[2272]  = 1;
  ram[2273]  = 1;
  ram[2274]  = 1;
  ram[2275]  = 1;
  ram[2276]  = 1;
  ram[2277]  = 1;
  ram[2278]  = 1;
  ram[2279]  = 1;
  ram[2280]  = 1;
  ram[2281]  = 1;
  ram[2282]  = 1;
  ram[2283]  = 1;
  ram[2284]  = 1;
  ram[2285]  = 1;
  ram[2286]  = 1;
  ram[2287]  = 1;
  ram[2288]  = 1;
  ram[2289]  = 1;
  ram[2290]  = 1;
  ram[2291]  = 1;
  ram[2292]  = 1;
  ram[2293]  = 1;
  ram[2294]  = 1;
  ram[2295]  = 1;
  ram[2296]  = 1;
  ram[2297]  = 1;
  ram[2298]  = 1;
  ram[2299]  = 1;
  ram[2300]  = 1;
  ram[2301]  = 1;
  ram[2302]  = 1;
  ram[2303]  = 1;
  ram[2304]  = 1;
  ram[2305]  = 1;
  ram[2306]  = 1;
  ram[2307]  = 1;
  ram[2308]  = 1;
  ram[2309]  = 1;
  ram[2310]  = 1;
  ram[2311]  = 1;
  ram[2312]  = 1;
  ram[2313]  = 1;
  ram[2314]  = 1;
  ram[2315]  = 1;
  ram[2316]  = 1;
  ram[2317]  = 1;
  ram[2318]  = 1;
  ram[2319]  = 1;
  ram[2320]  = 1;
  ram[2321]  = 1;
  ram[2322]  = 1;
  ram[2323]  = 1;
  ram[2324]  = 1;
  ram[2325]  = 1;
  ram[2326]  = 1;
  ram[2327]  = 1;
  ram[2328]  = 1;
  ram[2329]  = 1;
  ram[2330]  = 1;
  ram[2331]  = 1;
  ram[2332]  = 1;
  ram[2333]  = 1;
  ram[2334]  = 1;
  ram[2335]  = 1;
  ram[2336]  = 1;
  ram[2337]  = 1;
  ram[2338]  = 1;
  ram[2339]  = 1;
  ram[2340]  = 1;
  ram[2341]  = 1;
  ram[2342]  = 1;
  ram[2343]  = 1;
  ram[2344]  = 1;
  ram[2345]  = 1;
  ram[2346]  = 1;
  ram[2347]  = 1;
  ram[2348]  = 1;
  ram[2349]  = 1;
  ram[2350]  = 1;
  ram[2351]  = 1;
  ram[2352]  = 1;
  ram[2353]  = 1;
  ram[2354]  = 1;
  ram[2355]  = 1;
  ram[2356]  = 1;
  ram[2357]  = 1;
  ram[2358]  = 1;
  ram[2359]  = 1;
  ram[2360]  = 1;
  ram[2361]  = 1;
  ram[2362]  = 1;
  ram[2363]  = 1;
  ram[2364]  = 1;
  ram[2365]  = 1;
  ram[2366]  = 1;
  ram[2367]  = 1;
  ram[2368]  = 1;
  ram[2369]  = 1;
  ram[2370]  = 1;
  ram[2371]  = 1;
  ram[2372]  = 1;
  ram[2373]  = 1;
  ram[2374]  = 1;
  ram[2375]  = 1;
  ram[2376]  = 1;
  ram[2377]  = 1;
  ram[2378]  = 1;
  ram[2379]  = 1;
  ram[2380]  = 1;
  ram[2381]  = 1;
  ram[2382]  = 1;
  ram[2383]  = 1;
  ram[2384]  = 1;
  ram[2385]  = 1;
  ram[2386]  = 1;
  ram[2387]  = 1;
  ram[2388]  = 1;
  ram[2389]  = 1;
  ram[2390]  = 1;
  ram[2391]  = 1;
  ram[2392]  = 1;
  ram[2393]  = 1;
  ram[2394]  = 1;
  ram[2395]  = 1;
  ram[2396]  = 1;
  ram[2397]  = 1;
  ram[2398]  = 1;
  ram[2399]  = 1;
  ram[2400]  = 1;
  ram[2401]  = 1;
  ram[2402]  = 1;
  ram[2403]  = 1;
  ram[2404]  = 1;
  ram[2405]  = 1;
  ram[2406]  = 1;
  ram[2407]  = 1;
  ram[2408]  = 1;
  ram[2409]  = 1;
  ram[2410]  = 1;
  ram[2411]  = 1;
  ram[2412]  = 1;
  ram[2413]  = 1;
  ram[2414]  = 1;
  ram[2415]  = 1;
  ram[2416]  = 1;
  ram[2417]  = 1;
  ram[2418]  = 1;
  ram[2419]  = 1;
  ram[2420]  = 1;
  ram[2421]  = 1;
  ram[2422]  = 1;
  ram[2423]  = 1;
  ram[2424]  = 1;
  ram[2425]  = 1;
  ram[2426]  = 1;
  ram[2427]  = 1;
  ram[2428]  = 1;
  ram[2429]  = 1;
  ram[2430]  = 1;
  ram[2431]  = 1;
  ram[2432]  = 1;
  ram[2433]  = 1;
  ram[2434]  = 1;
  ram[2435]  = 1;
  ram[2436]  = 1;
  ram[2437]  = 1;
  ram[2438]  = 1;
  ram[2439]  = 1;
  ram[2440]  = 1;
  ram[2441]  = 1;
  ram[2442]  = 1;
  ram[2443]  = 1;
  ram[2444]  = 1;
  ram[2445]  = 1;
  ram[2446]  = 1;
  ram[2447]  = 1;
  ram[2448]  = 1;
  ram[2449]  = 1;
  ram[2450]  = 1;
  ram[2451]  = 1;
  ram[2452]  = 1;
  ram[2453]  = 1;
  ram[2454]  = 1;
  ram[2455]  = 1;
  ram[2456]  = 1;
  ram[2457]  = 1;
  ram[2458]  = 1;
  ram[2459]  = 1;
  ram[2460]  = 1;
  ram[2461]  = 1;
  ram[2462]  = 1;
  ram[2463]  = 1;
  ram[2464]  = 1;
  ram[2465]  = 1;
  ram[2466]  = 1;
  ram[2467]  = 1;
  ram[2468]  = 1;
  ram[2469]  = 1;
  ram[2470]  = 1;
  ram[2471]  = 1;
  ram[2472]  = 1;
  ram[2473]  = 1;
  ram[2474]  = 1;
  ram[2475]  = 1;
  ram[2476]  = 1;
  ram[2477]  = 1;
  ram[2478]  = 1;
  ram[2479]  = 1;
  ram[2480]  = 1;
  ram[2481]  = 1;
  ram[2482]  = 1;
  ram[2483]  = 1;
  ram[2484]  = 1;
  ram[2485]  = 1;
  ram[2486]  = 1;
  ram[2487]  = 1;
  ram[2488]  = 1;
  ram[2489]  = 1;
  ram[2490]  = 1;
  ram[2491]  = 1;
  ram[2492]  = 1;
  ram[2493]  = 1;
  ram[2494]  = 1;
  ram[2495]  = 1;
  ram[2496]  = 1;
  ram[2497]  = 1;
  ram[2498]  = 1;
  ram[2499]  = 1;
  ram[2500]  = 1;
  ram[2501]  = 1;
  ram[2502]  = 1;
  ram[2503]  = 1;
  ram[2504]  = 1;
  ram[2505]  = 1;
  ram[2506]  = 1;
  ram[2507]  = 1;
  ram[2508]  = 1;
  ram[2509]  = 1;
  ram[2510]  = 1;
  ram[2511]  = 1;
  ram[2512]  = 1;
  ram[2513]  = 1;
  ram[2514]  = 1;
  ram[2515]  = 1;
  ram[2516]  = 1;
  ram[2517]  = 1;
  ram[2518]  = 1;
  ram[2519]  = 1;
  ram[2520]  = 1;
  ram[2521]  = 1;
  ram[2522]  = 1;
  ram[2523]  = 1;
  ram[2524]  = 1;
  ram[2525]  = 1;
  ram[2526]  = 1;
  ram[2527]  = 1;
  ram[2528]  = 1;
  ram[2529]  = 1;
  ram[2530]  = 1;
  ram[2531]  = 1;
  ram[2532]  = 1;
  ram[2533]  = 1;
  ram[2534]  = 1;
  ram[2535]  = 1;
  ram[2536]  = 1;
  ram[2537]  = 1;
  ram[2538]  = 1;
  ram[2539]  = 1;
  ram[2540]  = 1;
  ram[2541]  = 1;
  ram[2542]  = 1;
  ram[2543]  = 1;
  ram[2544]  = 1;
  ram[2545]  = 1;
  ram[2546]  = 1;
  ram[2547]  = 1;
  ram[2548]  = 1;
  ram[2549]  = 1;
  ram[2550]  = 1;
  ram[2551]  = 1;
  ram[2552]  = 1;
  ram[2553]  = 1;
  ram[2554]  = 1;
  ram[2555]  = 1;
  ram[2556]  = 1;
  ram[2557]  = 1;
  ram[2558]  = 1;
  ram[2559]  = 1;
  ram[2560]  = 1;
  ram[2561]  = 1;
  ram[2562]  = 1;
  ram[2563]  = 1;
  ram[2564]  = 1;
  ram[2565]  = 1;
  ram[2566]  = 1;
  ram[2567]  = 1;
  ram[2568]  = 1;
  ram[2569]  = 1;
  ram[2570]  = 1;
  ram[2571]  = 1;
  ram[2572]  = 1;
  ram[2573]  = 1;
  ram[2574]  = 1;
  ram[2575]  = 1;
  ram[2576]  = 1;
  ram[2577]  = 1;
  ram[2578]  = 1;
  ram[2579]  = 1;
  ram[2580]  = 1;
  ram[2581]  = 1;
  ram[2582]  = 1;
  ram[2583]  = 1;
  ram[2584]  = 1;
  ram[2585]  = 1;
  ram[2586]  = 1;
  ram[2587]  = 1;
  ram[2588]  = 1;
  ram[2589]  = 1;
  ram[2590]  = 1;
  ram[2591]  = 1;
  ram[2592]  = 1;
  ram[2593]  = 1;
  ram[2594]  = 1;
  ram[2595]  = 1;
  ram[2596]  = 1;
  ram[2597]  = 1;
  ram[2598]  = 1;
  ram[2599]  = 1;
  ram[2600]  = 1;
  ram[2601]  = 1;
  ram[2602]  = 1;
  ram[2603]  = 1;
  ram[2604]  = 1;
  ram[2605]  = 1;
  ram[2606]  = 1;
  ram[2607]  = 1;
  ram[2608]  = 1;
  ram[2609]  = 1;
  ram[2610]  = 1;
  ram[2611]  = 1;
  ram[2612]  = 1;
  ram[2613]  = 1;
  ram[2614]  = 1;
  ram[2615]  = 1;
  ram[2616]  = 1;
  ram[2617]  = 1;
  ram[2618]  = 1;
  ram[2619]  = 1;
  ram[2620]  = 1;
  ram[2621]  = 1;
  ram[2622]  = 1;
  ram[2623]  = 1;
  ram[2624]  = 1;
  ram[2625]  = 1;
  ram[2626]  = 1;
  ram[2627]  = 1;
  ram[2628]  = 1;
  ram[2629]  = 1;
  ram[2630]  = 1;
  ram[2631]  = 1;
  ram[2632]  = 1;
  ram[2633]  = 1;
  ram[2634]  = 1;
  ram[2635]  = 1;
  ram[2636]  = 1;
  ram[2637]  = 1;
  ram[2638]  = 1;
  ram[2639]  = 1;
  ram[2640]  = 1;
  ram[2641]  = 1;
  ram[2642]  = 1;
  ram[2643]  = 1;
  ram[2644]  = 1;
  ram[2645]  = 1;
  ram[2646]  = 1;
  ram[2647]  = 1;
  ram[2648]  = 1;
  ram[2649]  = 1;
  ram[2650]  = 1;
  ram[2651]  = 1;
  ram[2652]  = 1;
  ram[2653]  = 1;
  ram[2654]  = 1;
  ram[2655]  = 1;
  ram[2656]  = 1;
  ram[2657]  = 1;
  ram[2658]  = 1;
  ram[2659]  = 1;
  ram[2660]  = 1;
  ram[2661]  = 1;
  ram[2662]  = 1;
  ram[2663]  = 1;
  ram[2664]  = 1;
  ram[2665]  = 1;
  ram[2666]  = 1;
  ram[2667]  = 1;
  ram[2668]  = 1;
  ram[2669]  = 1;
  ram[2670]  = 1;
  ram[2671]  = 1;
  ram[2672]  = 1;
  ram[2673]  = 1;
  ram[2674]  = 1;
  ram[2675]  = 1;
  ram[2676]  = 1;
  ram[2677]  = 1;
  ram[2678]  = 1;
  ram[2679]  = 1;
  ram[2680]  = 1;
  ram[2681]  = 1;
  ram[2682]  = 1;
  ram[2683]  = 1;
  ram[2684]  = 1;
  ram[2685]  = 1;
  ram[2686]  = 1;
  ram[2687]  = 1;
  ram[2688]  = 1;
  ram[2689]  = 1;
  ram[2690]  = 1;
  ram[2691]  = 1;
  ram[2692]  = 1;
  ram[2693]  = 1;
  ram[2694]  = 1;
  ram[2695]  = 1;
  ram[2696]  = 1;
  ram[2697]  = 1;
  ram[2698]  = 1;
  ram[2699]  = 1;
  ram[2700]  = 1;
  ram[2701]  = 1;
  ram[2702]  = 1;
  ram[2703]  = 1;
  ram[2704]  = 1;
  ram[2705]  = 1;
  ram[2706]  = 1;
  ram[2707]  = 1;
  ram[2708]  = 1;
  ram[2709]  = 1;
  ram[2710]  = 1;
  ram[2711]  = 1;
  ram[2712]  = 1;
  ram[2713]  = 1;
  ram[2714]  = 1;
  ram[2715]  = 1;
  ram[2716]  = 1;
  ram[2717]  = 1;
  ram[2718]  = 1;
  ram[2719]  = 1;
  ram[2720]  = 1;
  ram[2721]  = 1;
  ram[2722]  = 1;
  ram[2723]  = 1;
  ram[2724]  = 1;
  ram[2725]  = 1;
  ram[2726]  = 1;
  ram[2727]  = 1;
  ram[2728]  = 1;
  ram[2729]  = 1;
  ram[2730]  = 1;
  ram[2731]  = 1;
  ram[2732]  = 1;
  ram[2733]  = 1;
  ram[2734]  = 1;
  ram[2735]  = 1;
  ram[2736]  = 1;
  ram[2737]  = 1;
  ram[2738]  = 1;
  ram[2739]  = 1;
  ram[2740]  = 1;
  ram[2741]  = 1;
  ram[2742]  = 1;
  ram[2743]  = 1;
  ram[2744]  = 1;
  ram[2745]  = 1;
  ram[2746]  = 1;
  ram[2747]  = 1;
  ram[2748]  = 1;
  ram[2749]  = 1;
  ram[2750]  = 1;
  ram[2751]  = 1;
  ram[2752]  = 1;
  ram[2753]  = 1;
  ram[2754]  = 1;
  ram[2755]  = 1;
  ram[2756]  = 1;
  ram[2757]  = 1;
  ram[2758]  = 1;
  ram[2759]  = 1;
  ram[2760]  = 1;
  ram[2761]  = 1;
  ram[2762]  = 1;
  ram[2763]  = 1;
  ram[2764]  = 1;
  ram[2765]  = 1;
  ram[2766]  = 1;
  ram[2767]  = 1;
  ram[2768]  = 1;
  ram[2769]  = 1;
  ram[2770]  = 1;
  ram[2771]  = 1;
  ram[2772]  = 1;
  ram[2773]  = 1;
  ram[2774]  = 1;
  ram[2775]  = 1;
  ram[2776]  = 1;
  ram[2777]  = 1;
  ram[2778]  = 1;
  ram[2779]  = 1;
  ram[2780]  = 1;
  ram[2781]  = 1;
  ram[2782]  = 1;
  ram[2783]  = 1;
  ram[2784]  = 1;
  ram[2785]  = 1;
  ram[2786]  = 1;
  ram[2787]  = 1;
  ram[2788]  = 1;
  ram[2789]  = 1;
  ram[2790]  = 1;
  ram[2791]  = 1;
  ram[2792]  = 1;
  ram[2793]  = 1;
  ram[2794]  = 1;
  ram[2795]  = 1;
  ram[2796]  = 1;
  ram[2797]  = 1;
  ram[2798]  = 1;
  ram[2799]  = 1;
  ram[2800]  = 1;
  ram[2801]  = 1;
  ram[2802]  = 1;
  ram[2803]  = 1;
  ram[2804]  = 1;
  ram[2805]  = 1;
  ram[2806]  = 1;
  ram[2807]  = 1;
  ram[2808]  = 1;
  ram[2809]  = 1;
  ram[2810]  = 1;
  ram[2811]  = 1;
  ram[2812]  = 1;
  ram[2813]  = 1;
  ram[2814]  = 1;
  ram[2815]  = 1;
  ram[2816]  = 1;
  ram[2817]  = 1;
  ram[2818]  = 1;
  ram[2819]  = 1;
  ram[2820]  = 1;
  ram[2821]  = 1;
  ram[2822]  = 1;
  ram[2823]  = 1;
  ram[2824]  = 1;
  ram[2825]  = 1;
  ram[2826]  = 1;
  ram[2827]  = 1;
  ram[2828]  = 1;
  ram[2829]  = 1;
  ram[2830]  = 1;
  ram[2831]  = 1;
  ram[2832]  = 1;
  ram[2833]  = 1;
  ram[2834]  = 1;
  ram[2835]  = 1;
  ram[2836]  = 1;
  ram[2837]  = 1;
  ram[2838]  = 1;
  ram[2839]  = 1;
  ram[2840]  = 1;
  ram[2841]  = 1;
  ram[2842]  = 1;
  ram[2843]  = 1;
  ram[2844]  = 1;
  ram[2845]  = 1;
  ram[2846]  = 1;
  ram[2847]  = 1;
  ram[2848]  = 1;
  ram[2849]  = 1;
  ram[2850]  = 1;
  ram[2851]  = 1;
  ram[2852]  = 1;
  ram[2853]  = 1;
  ram[2854]  = 1;
  ram[2855]  = 1;
  ram[2856]  = 1;
  ram[2857]  = 1;
  ram[2858]  = 1;
  ram[2859]  = 1;
  ram[2860]  = 1;
  ram[2861]  = 1;
  ram[2862]  = 1;
  ram[2863]  = 1;
  ram[2864]  = 1;
  ram[2865]  = 1;
  ram[2866]  = 1;
  ram[2867]  = 1;
  ram[2868]  = 1;
  ram[2869]  = 1;
  ram[2870]  = 1;
  ram[2871]  = 1;
  ram[2872]  = 1;
  ram[2873]  = 1;
  ram[2874]  = 1;
  ram[2875]  = 1;
  ram[2876]  = 1;
  ram[2877]  = 1;
  ram[2878]  = 1;
  ram[2879]  = 1;
  ram[2880]  = 1;
  ram[2881]  = 1;
  ram[2882]  = 1;
  ram[2883]  = 1;
  ram[2884]  = 1;
  ram[2885]  = 1;
  ram[2886]  = 1;
  ram[2887]  = 1;
  ram[2888]  = 1;
  ram[2889]  = 1;
  ram[2890]  = 1;
  ram[2891]  = 1;
  ram[2892]  = 1;
  ram[2893]  = 1;
  ram[2894]  = 1;
  ram[2895]  = 1;
  ram[2896]  = 1;
  ram[2897]  = 1;
  ram[2898]  = 1;
  ram[2899]  = 1;
  ram[2900]  = 1;
  ram[2901]  = 1;
  ram[2902]  = 1;
  ram[2903]  = 1;
  ram[2904]  = 1;
  ram[2905]  = 1;
  ram[2906]  = 1;
  ram[2907]  = 1;
  ram[2908]  = 1;
  ram[2909]  = 1;
  ram[2910]  = 1;
  ram[2911]  = 1;
  ram[2912]  = 1;
  ram[2913]  = 1;
  ram[2914]  = 1;
  ram[2915]  = 1;
  ram[2916]  = 1;
  ram[2917]  = 1;
  ram[2918]  = 1;
  ram[2919]  = 1;
  ram[2920]  = 1;
  ram[2921]  = 1;
  ram[2922]  = 1;
  ram[2923]  = 1;
  ram[2924]  = 1;
  ram[2925]  = 1;
  ram[2926]  = 1;
  ram[2927]  = 1;
  ram[2928]  = 1;
  ram[2929]  = 1;
  ram[2930]  = 1;
  ram[2931]  = 1;
  ram[2932]  = 1;
  ram[2933]  = 1;
  ram[2934]  = 1;
  ram[2935]  = 1;
  ram[2936]  = 1;
  ram[2937]  = 1;
  ram[2938]  = 1;
  ram[2939]  = 1;
  ram[2940]  = 1;
  ram[2941]  = 1;
  ram[2942]  = 1;
  ram[2943]  = 1;
  ram[2944]  = 1;
  ram[2945]  = 1;
  ram[2946]  = 1;
  ram[2947]  = 1;
  ram[2948]  = 1;
  ram[2949]  = 1;
  ram[2950]  = 1;
  ram[2951]  = 1;
  ram[2952]  = 1;
  ram[2953]  = 1;
  ram[2954]  = 1;
  ram[2955]  = 1;
  ram[2956]  = 1;
  ram[2957]  = 1;
  ram[2958]  = 1;
  ram[2959]  = 1;
  ram[2960]  = 1;
  ram[2961]  = 1;
  ram[2962]  = 1;
  ram[2963]  = 1;
  ram[2964]  = 1;
  ram[2965]  = 1;
  ram[2966]  = 1;
  ram[2967]  = 1;
  ram[2968]  = 1;
  ram[2969]  = 1;
  ram[2970]  = 1;
  ram[2971]  = 1;
  ram[2972]  = 1;
  ram[2973]  = 1;
  ram[2974]  = 1;
  ram[2975]  = 1;
  ram[2976]  = 1;
  ram[2977]  = 1;
  ram[2978]  = 1;
  ram[2979]  = 1;
  ram[2980]  = 1;
  ram[2981]  = 1;
  ram[2982]  = 1;
  ram[2983]  = 1;
  ram[2984]  = 1;
  ram[2985]  = 1;
  ram[2986]  = 1;
  ram[2987]  = 1;
  ram[2988]  = 1;
  ram[2989]  = 1;
  ram[2990]  = 1;
  ram[2991]  = 1;
  ram[2992]  = 1;
  ram[2993]  = 1;
  ram[2994]  = 1;
  ram[2995]  = 1;
  ram[2996]  = 1;
  ram[2997]  = 1;
  ram[2998]  = 1;
  ram[2999]  = 1;
  ram[3000]  = 1;
  ram[3001]  = 1;
  ram[3002]  = 1;
  ram[3003]  = 1;
  ram[3004]  = 1;
  ram[3005]  = 1;
  ram[3006]  = 1;
  ram[3007]  = 1;
  ram[3008]  = 1;
  ram[3009]  = 1;
  ram[3010]  = 1;
  ram[3011]  = 1;
  ram[3012]  = 1;
  ram[3013]  = 1;
  ram[3014]  = 1;
  ram[3015]  = 1;
  ram[3016]  = 1;
  ram[3017]  = 1;
  ram[3018]  = 1;
  ram[3019]  = 1;
  ram[3020]  = 1;
  ram[3021]  = 1;
  ram[3022]  = 1;
  ram[3023]  = 1;
  ram[3024]  = 1;
  ram[3025]  = 1;
  ram[3026]  = 1;
  ram[3027]  = 1;
  ram[3028]  = 1;
  ram[3029]  = 1;
  ram[3030]  = 1;
  ram[3031]  = 1;
  ram[3032]  = 1;
  ram[3033]  = 1;
  ram[3034]  = 1;
  ram[3035]  = 1;
  ram[3036]  = 1;
  ram[3037]  = 1;
  ram[3038]  = 1;
  ram[3039]  = 1;
  ram[3040]  = 1;
  ram[3041]  = 1;
  ram[3042]  = 1;
  ram[3043]  = 1;
  ram[3044]  = 1;
  ram[3045]  = 1;
  ram[3046]  = 1;
  ram[3047]  = 1;
  ram[3048]  = 1;
  ram[3049]  = 1;
  ram[3050]  = 1;
  ram[3051]  = 1;
  ram[3052]  = 1;
  ram[3053]  = 1;
  ram[3054]  = 1;
  ram[3055]  = 1;
  ram[3056]  = 1;
  ram[3057]  = 1;
  ram[3058]  = 1;
  ram[3059]  = 1;
  ram[3060]  = 1;
  ram[3061]  = 1;
  ram[3062]  = 1;
  ram[3063]  = 1;
  ram[3064]  = 1;
  ram[3065]  = 1;
  ram[3066]  = 1;
  ram[3067]  = 1;
  ram[3068]  = 1;
  ram[3069]  = 1;
  ram[3070]  = 1;
  ram[3071]  = 1;
  ram[3072]  = 1;
  ram[3073]  = 1;
  ram[3074]  = 1;
  ram[3075]  = 1;
  ram[3076]  = 1;
  ram[3077]  = 1;
  ram[3078]  = 1;
  ram[3079]  = 1;
  ram[3080]  = 1;
  ram[3081]  = 1;
  ram[3082]  = 1;
  ram[3083]  = 1;
  ram[3084]  = 1;
  ram[3085]  = 1;
  ram[3086]  = 1;
  ram[3087]  = 1;
  ram[3088]  = 1;
  ram[3089]  = 1;
  ram[3090]  = 1;
  ram[3091]  = 1;
  ram[3092]  = 1;
  ram[3093]  = 1;
  ram[3094]  = 1;
  ram[3095]  = 1;
  ram[3096]  = 1;
  ram[3097]  = 1;
  ram[3098]  = 1;
  ram[3099]  = 1;
  ram[3100]  = 1;
  ram[3101]  = 1;
  ram[3102]  = 1;
  ram[3103]  = 1;
  ram[3104]  = 1;
  ram[3105]  = 1;
  ram[3106]  = 1;
  ram[3107]  = 1;
  ram[3108]  = 1;
  ram[3109]  = 1;
  ram[3110]  = 1;
  ram[3111]  = 1;
  ram[3112]  = 1;
  ram[3113]  = 1;
  ram[3114]  = 1;
  ram[3115]  = 1;
  ram[3116]  = 1;
  ram[3117]  = 1;
  ram[3118]  = 1;
  ram[3119]  = 1;
  ram[3120]  = 1;
  ram[3121]  = 1;
  ram[3122]  = 1;
  ram[3123]  = 1;
  ram[3124]  = 1;
  ram[3125]  = 1;
  ram[3126]  = 1;
  ram[3127]  = 1;
  ram[3128]  = 1;
  ram[3129]  = 1;
  ram[3130]  = 1;
  ram[3131]  = 1;
  ram[3132]  = 1;
  ram[3133]  = 1;
  ram[3134]  = 1;
  ram[3135]  = 1;
  ram[3136]  = 1;
  ram[3137]  = 1;
  ram[3138]  = 1;
  ram[3139]  = 1;
  ram[3140]  = 1;
  ram[3141]  = 1;
  ram[3142]  = 1;
  ram[3143]  = 1;
  ram[3144]  = 1;
  ram[3145]  = 1;
  ram[3146]  = 1;
  ram[3147]  = 1;
  ram[3148]  = 1;
  ram[3149]  = 1;
  ram[3150]  = 1;
  ram[3151]  = 1;
  ram[3152]  = 1;
  ram[3153]  = 1;
  ram[3154]  = 1;
  ram[3155]  = 1;
  ram[3156]  = 1;
  ram[3157]  = 1;
  ram[3158]  = 1;
  ram[3159]  = 1;
  ram[3160]  = 1;
  ram[3161]  = 1;
  ram[3162]  = 1;
  ram[3163]  = 1;
  ram[3164]  = 1;
  ram[3165]  = 1;
  ram[3166]  = 1;
  ram[3167]  = 1;
  ram[3168]  = 1;
  ram[3169]  = 1;
  ram[3170]  = 1;
  ram[3171]  = 1;
  ram[3172]  = 1;
  ram[3173]  = 1;
  ram[3174]  = 1;
  ram[3175]  = 1;
  ram[3176]  = 1;
  ram[3177]  = 1;
  ram[3178]  = 1;
  ram[3179]  = 1;
  ram[3180]  = 1;
  ram[3181]  = 1;
  ram[3182]  = 1;
  ram[3183]  = 1;
  ram[3184]  = 1;
  ram[3185]  = 1;
  ram[3186]  = 1;
  ram[3187]  = 1;
  ram[3188]  = 1;
  ram[3189]  = 1;
  ram[3190]  = 1;
  ram[3191]  = 1;
  ram[3192]  = 1;
  ram[3193]  = 1;
  ram[3194]  = 1;
  ram[3195]  = 1;
  ram[3196]  = 1;
  ram[3197]  = 1;
  ram[3198]  = 1;
  ram[3199]  = 1;
  ram[3200]  = 1;
  ram[3201]  = 1;
  ram[3202]  = 1;
  ram[3203]  = 1;
  ram[3204]  = 1;
  ram[3205]  = 1;
  ram[3206]  = 1;
  ram[3207]  = 1;
  ram[3208]  = 1;
  ram[3209]  = 1;
  ram[3210]  = 1;
  ram[3211]  = 1;
  ram[3212]  = 1;
  ram[3213]  = 1;
  ram[3214]  = 1;
  ram[3215]  = 1;
  ram[3216]  = 1;
  ram[3217]  = 1;
  ram[3218]  = 1;
  ram[3219]  = 1;
  ram[3220]  = 1;
  ram[3221]  = 1;
  ram[3222]  = 1;
  ram[3223]  = 1;
  ram[3224]  = 1;
  ram[3225]  = 1;
  ram[3226]  = 1;
  ram[3227]  = 1;
  ram[3228]  = 1;
  ram[3229]  = 1;
  ram[3230]  = 1;
  ram[3231]  = 1;
  ram[3232]  = 1;
  ram[3233]  = 1;
  ram[3234]  = 1;
  ram[3235]  = 1;
  ram[3236]  = 1;
  ram[3237]  = 1;
  ram[3238]  = 1;
  ram[3239]  = 1;
  ram[3240]  = 1;
  ram[3241]  = 1;
  ram[3242]  = 1;
  ram[3243]  = 1;
  ram[3244]  = 1;
  ram[3245]  = 1;
  ram[3246]  = 1;
  ram[3247]  = 1;
  ram[3248]  = 1;
  ram[3249]  = 1;
  ram[3250]  = 1;
  ram[3251]  = 1;
  ram[3252]  = 1;
  ram[3253]  = 1;
  ram[3254]  = 1;
  ram[3255]  = 1;
  ram[3256]  = 1;
  ram[3257]  = 1;
  ram[3258]  = 1;
  ram[3259]  = 1;
  ram[3260]  = 1;
  ram[3261]  = 1;
  ram[3262]  = 1;
  ram[3263]  = 1;
  ram[3264]  = 1;
  ram[3265]  = 1;
  ram[3266]  = 1;
  ram[3267]  = 1;
  ram[3268]  = 1;
  ram[3269]  = 1;
  ram[3270]  = 1;
  ram[3271]  = 1;
  ram[3272]  = 1;
  ram[3273]  = 1;
  ram[3274]  = 1;
  ram[3275]  = 1;
  ram[3276]  = 1;
  ram[3277]  = 1;
  ram[3278]  = 1;
  ram[3279]  = 1;
  ram[3280]  = 1;
  ram[3281]  = 1;
  ram[3282]  = 1;
  ram[3283]  = 1;
  ram[3284]  = 1;
  ram[3285]  = 1;
  ram[3286]  = 1;
  ram[3287]  = 1;
  ram[3288]  = 1;
  ram[3289]  = 1;
  ram[3290]  = 1;
  ram[3291]  = 1;
  ram[3292]  = 1;
  ram[3293]  = 1;
  ram[3294]  = 1;
  ram[3295]  = 1;
  ram[3296]  = 1;
  ram[3297]  = 1;
  ram[3298]  = 1;
  ram[3299]  = 1;
  ram[3300]  = 1;
  ram[3301]  = 1;
  ram[3302]  = 1;
  ram[3303]  = 1;
  ram[3304]  = 1;
  ram[3305]  = 1;
  ram[3306]  = 1;
  ram[3307]  = 1;
  ram[3308]  = 1;
  ram[3309]  = 1;
  ram[3310]  = 1;
  ram[3311]  = 1;
  ram[3312]  = 1;
  ram[3313]  = 1;
  ram[3314]  = 1;
  ram[3315]  = 1;
  ram[3316]  = 1;
  ram[3317]  = 1;
  ram[3318]  = 1;
  ram[3319]  = 1;
  ram[3320]  = 1;
  ram[3321]  = 1;
  ram[3322]  = 1;
  ram[3323]  = 1;
  ram[3324]  = 1;
  ram[3325]  = 1;
  ram[3326]  = 1;
  ram[3327]  = 1;
  ram[3328]  = 1;
  ram[3329]  = 1;
  ram[3330]  = 1;
  ram[3331]  = 1;
  ram[3332]  = 1;
  ram[3333]  = 1;
  ram[3334]  = 1;
  ram[3335]  = 1;
  ram[3336]  = 1;
  ram[3337]  = 1;
  ram[3338]  = 1;
  ram[3339]  = 1;
  ram[3340]  = 1;
  ram[3341]  = 1;
  ram[3342]  = 1;
  ram[3343]  = 1;
  ram[3344]  = 1;
  ram[3345]  = 1;
  ram[3346]  = 1;
  ram[3347]  = 1;
  ram[3348]  = 1;
  ram[3349]  = 1;
  ram[3350]  = 1;
  ram[3351]  = 1;
  ram[3352]  = 1;
  ram[3353]  = 1;
  ram[3354]  = 1;
  ram[3355]  = 1;
  ram[3356]  = 1;
  ram[3357]  = 1;
  ram[3358]  = 1;
  ram[3359]  = 1;
  ram[3360]  = 1;
  ram[3361]  = 1;
  ram[3362]  = 1;
  ram[3363]  = 1;
  ram[3364]  = 1;
  ram[3365]  = 1;
  ram[3366]  = 1;
  ram[3367]  = 1;
  ram[3368]  = 1;
  ram[3369]  = 1;
  ram[3370]  = 1;
  ram[3371]  = 1;
  ram[3372]  = 1;
  ram[3373]  = 1;
  ram[3374]  = 1;
  ram[3375]  = 1;
  ram[3376]  = 1;
  ram[3377]  = 1;
  ram[3378]  = 1;
  ram[3379]  = 1;
  ram[3380]  = 1;
  ram[3381]  = 1;
  ram[3382]  = 1;
  ram[3383]  = 1;
  ram[3384]  = 1;
  ram[3385]  = 1;
  ram[3386]  = 1;
  ram[3387]  = 1;
  ram[3388]  = 1;
  ram[3389]  = 1;
  ram[3390]  = 1;
  ram[3391]  = 1;
  ram[3392]  = 1;
  ram[3393]  = 1;
  ram[3394]  = 1;
  ram[3395]  = 1;
  ram[3396]  = 1;
  ram[3397]  = 1;
  ram[3398]  = 1;
  ram[3399]  = 1;
  ram[3400]  = 1;
  ram[3401]  = 1;
  ram[3402]  = 1;
  ram[3403]  = 1;
  ram[3404]  = 1;
  ram[3405]  = 1;
  ram[3406]  = 1;
  ram[3407]  = 1;
  ram[3408]  = 1;
  ram[3409]  = 1;
  ram[3410]  = 1;
  ram[3411]  = 1;
  ram[3412]  = 1;
  ram[3413]  = 1;
  ram[3414]  = 1;
  ram[3415]  = 1;
  ram[3416]  = 1;
  ram[3417]  = 1;
  ram[3418]  = 1;
  ram[3419]  = 1;
  ram[3420]  = 1;
  ram[3421]  = 1;
  ram[3422]  = 1;
  ram[3423]  = 1;
  ram[3424]  = 1;
  ram[3425]  = 1;
  ram[3426]  = 1;
  ram[3427]  = 1;
  ram[3428]  = 1;
  ram[3429]  = 1;
  ram[3430]  = 1;
  ram[3431]  = 1;
  ram[3432]  = 1;
  ram[3433]  = 1;
  ram[3434]  = 1;
  ram[3435]  = 1;
  ram[3436]  = 1;
  ram[3437]  = 1;
  ram[3438]  = 1;
  ram[3439]  = 1;
  ram[3440]  = 1;
  ram[3441]  = 1;
  ram[3442]  = 1;
  ram[3443]  = 1;
  ram[3444]  = 1;
  ram[3445]  = 1;
  ram[3446]  = 1;
  ram[3447]  = 1;
  ram[3448]  = 1;
  ram[3449]  = 1;
  ram[3450]  = 1;
  ram[3451]  = 1;
  ram[3452]  = 1;
  ram[3453]  = 1;
  ram[3454]  = 1;
  ram[3455]  = 1;
  ram[3456]  = 1;
  ram[3457]  = 1;
  ram[3458]  = 1;
  ram[3459]  = 1;
  ram[3460]  = 1;
  ram[3461]  = 1;
  ram[3462]  = 1;
  ram[3463]  = 1;
  ram[3464]  = 1;
  ram[3465]  = 1;
  ram[3466]  = 1;
  ram[3467]  = 1;
  ram[3468]  = 1;
  ram[3469]  = 1;
  ram[3470]  = 1;
  ram[3471]  = 1;
  ram[3472]  = 1;
  ram[3473]  = 1;
  ram[3474]  = 1;
  ram[3475]  = 1;
  ram[3476]  = 1;
  ram[3477]  = 1;
  ram[3478]  = 1;
  ram[3479]  = 1;
  ram[3480]  = 1;
  ram[3481]  = 1;
  ram[3482]  = 1;
  ram[3483]  = 1;
  ram[3484]  = 1;
  ram[3485]  = 1;
  ram[3486]  = 1;
  ram[3487]  = 1;
  ram[3488]  = 1;
  ram[3489]  = 1;
  ram[3490]  = 1;
  ram[3491]  = 1;
  ram[3492]  = 1;
  ram[3493]  = 1;
  ram[3494]  = 1;
  ram[3495]  = 1;
  ram[3496]  = 1;
  ram[3497]  = 1;
  ram[3498]  = 1;
  ram[3499]  = 1;
  ram[3500]  = 1;
  ram[3501]  = 1;
  ram[3502]  = 1;
  ram[3503]  = 1;
  ram[3504]  = 1;
  ram[3505]  = 1;
  ram[3506]  = 1;
  ram[3507]  = 1;
  ram[3508]  = 1;
  ram[3509]  = 1;
  ram[3510]  = 1;
  ram[3511]  = 1;
  ram[3512]  = 1;
  ram[3513]  = 1;
  ram[3514]  = 1;
  ram[3515]  = 1;
  ram[3516]  = 1;
  ram[3517]  = 1;
  ram[3518]  = 1;
  ram[3519]  = 1;
  ram[3520]  = 1;
  ram[3521]  = 1;
  ram[3522]  = 1;
  ram[3523]  = 1;
  ram[3524]  = 1;
  ram[3525]  = 1;
  ram[3526]  = 1;
  ram[3527]  = 1;
  ram[3528]  = 1;
  ram[3529]  = 1;
  ram[3530]  = 1;
  ram[3531]  = 1;
  ram[3532]  = 1;
  ram[3533]  = 1;
  ram[3534]  = 1;
  ram[3535]  = 1;
  ram[3536]  = 1;
  ram[3537]  = 1;
  ram[3538]  = 1;
  ram[3539]  = 1;
  ram[3540]  = 1;
  ram[3541]  = 1;
  ram[3542]  = 1;
  ram[3543]  = 1;
  ram[3544]  = 1;
  ram[3545]  = 1;
  ram[3546]  = 1;
  ram[3547]  = 1;
  ram[3548]  = 1;
  ram[3549]  = 1;
  ram[3550]  = 1;
  ram[3551]  = 1;
  ram[3552]  = 1;
  ram[3553]  = 1;
  ram[3554]  = 1;
  ram[3555]  = 1;
  ram[3556]  = 1;
  ram[3557]  = 1;
  ram[3558]  = 1;
  ram[3559]  = 1;
  ram[3560]  = 1;
  ram[3561]  = 1;
  ram[3562]  = 1;
  ram[3563]  = 1;
  ram[3564]  = 1;
  ram[3565]  = 1;
  ram[3566]  = 1;
  ram[3567]  = 1;
  ram[3568]  = 1;
  ram[3569]  = 1;
  ram[3570]  = 1;
  ram[3571]  = 1;
  ram[3572]  = 1;
  ram[3573]  = 1;
  ram[3574]  = 1;
  ram[3575]  = 1;
  ram[3576]  = 1;
  ram[3577]  = 1;
  ram[3578]  = 1;
  ram[3579]  = 1;
  ram[3580]  = 1;
  ram[3581]  = 1;
  ram[3582]  = 1;
  ram[3583]  = 1;
  ram[3584]  = 1;
  ram[3585]  = 1;
  ram[3586]  = 1;
  ram[3587]  = 1;
  ram[3588]  = 1;
  ram[3589]  = 1;
  ram[3590]  = 1;
  ram[3591]  = 1;
  ram[3592]  = 1;
  ram[3593]  = 1;
  ram[3594]  = 1;
  ram[3595]  = 1;
  ram[3596]  = 1;
  ram[3597]  = 1;
  ram[3598]  = 1;
  ram[3599]  = 1;
  ram[3600]  = 1;
  ram[3601]  = 1;
  ram[3602]  = 1;
  ram[3603]  = 1;
  ram[3604]  = 1;
  ram[3605]  = 1;
  ram[3606]  = 1;
  ram[3607]  = 1;
  ram[3608]  = 1;
  ram[3609]  = 1;
  ram[3610]  = 1;
  ram[3611]  = 1;
  ram[3612]  = 1;
  ram[3613]  = 1;
  ram[3614]  = 1;
  ram[3615]  = 1;
  ram[3616]  = 1;
  ram[3617]  = 1;
  ram[3618]  = 1;
  ram[3619]  = 1;
  ram[3620]  = 1;
  ram[3621]  = 1;
  ram[3622]  = 1;
  ram[3623]  = 1;
  ram[3624]  = 1;
  ram[3625]  = 1;
  ram[3626]  = 1;
  ram[3627]  = 1;
  ram[3628]  = 1;
  ram[3629]  = 1;
  ram[3630]  = 1;
  ram[3631]  = 1;
  ram[3632]  = 1;
  ram[3633]  = 1;
  ram[3634]  = 1;
  ram[3635]  = 1;
  ram[3636]  = 1;
  ram[3637]  = 1;
  ram[3638]  = 1;
  ram[3639]  = 1;
  ram[3640]  = 1;
  ram[3641]  = 1;
  ram[3642]  = 1;
  ram[3643]  = 1;
  ram[3644]  = 1;
  ram[3645]  = 1;
  ram[3646]  = 1;
  ram[3647]  = 1;
  ram[3648]  = 1;
  ram[3649]  = 1;
  ram[3650]  = 1;
  ram[3651]  = 1;
  ram[3652]  = 1;
  ram[3653]  = 1;
  ram[3654]  = 1;
  ram[3655]  = 1;
  ram[3656]  = 1;
  ram[3657]  = 1;
  ram[3658]  = 1;
  ram[3659]  = 1;
  ram[3660]  = 1;
  ram[3661]  = 1;
  ram[3662]  = 1;
  ram[3663]  = 1;
  ram[3664]  = 1;
  ram[3665]  = 1;
  ram[3666]  = 1;
  ram[3667]  = 1;
  ram[3668]  = 1;
  ram[3669]  = 1;
  ram[3670]  = 1;
  ram[3671]  = 1;
  ram[3672]  = 1;
  ram[3673]  = 1;
  ram[3674]  = 1;
  ram[3675]  = 1;
  ram[3676]  = 1;
  ram[3677]  = 1;
  ram[3678]  = 1;
  ram[3679]  = 1;
  ram[3680]  = 1;
  ram[3681]  = 1;
  ram[3682]  = 1;
  ram[3683]  = 1;
  ram[3684]  = 1;
  ram[3685]  = 1;
  ram[3686]  = 1;
  ram[3687]  = 1;
  ram[3688]  = 1;
  ram[3689]  = 1;
  ram[3690]  = 1;
  ram[3691]  = 1;
  ram[3692]  = 1;
  ram[3693]  = 1;
  ram[3694]  = 1;
  ram[3695]  = 1;
  ram[3696]  = 1;
  ram[3697]  = 1;
  ram[3698]  = 1;
  ram[3699]  = 1;
  ram[3700]  = 1;
  ram[3701]  = 1;
  ram[3702]  = 1;
  ram[3703]  = 1;
  ram[3704]  = 1;
  ram[3705]  = 1;
  ram[3706]  = 1;
  ram[3707]  = 1;
  ram[3708]  = 1;
  ram[3709]  = 1;
  ram[3710]  = 1;
  ram[3711]  = 1;
  ram[3712]  = 1;
  ram[3713]  = 1;
  ram[3714]  = 1;
  ram[3715]  = 1;
  ram[3716]  = 1;
  ram[3717]  = 1;
  ram[3718]  = 1;
  ram[3719]  = 1;
  ram[3720]  = 1;
  ram[3721]  = 1;
  ram[3722]  = 1;
  ram[3723]  = 1;
  ram[3724]  = 1;
  ram[3725]  = 1;
  ram[3726]  = 1;
  ram[3727]  = 1;
  ram[3728]  = 1;
  ram[3729]  = 1;
  ram[3730]  = 1;
  ram[3731]  = 1;
  ram[3732]  = 1;
  ram[3733]  = 1;
  ram[3734]  = 1;
  ram[3735]  = 1;
  ram[3736]  = 1;
  ram[3737]  = 1;
  ram[3738]  = 1;
  ram[3739]  = 1;
  ram[3740]  = 1;
  ram[3741]  = 1;
  ram[3742]  = 1;
  ram[3743]  = 1;
  ram[3744]  = 1;
  ram[3745]  = 1;
  ram[3746]  = 1;
  ram[3747]  = 1;
  ram[3748]  = 1;
  ram[3749]  = 1;
  ram[3750]  = 1;
  ram[3751]  = 1;
  ram[3752]  = 1;
  ram[3753]  = 1;
  ram[3754]  = 1;
  ram[3755]  = 1;
  ram[3756]  = 1;
  ram[3757]  = 1;
  ram[3758]  = 1;
  ram[3759]  = 1;
  ram[3760]  = 1;
  ram[3761]  = 1;
  ram[3762]  = 1;
  ram[3763]  = 1;
  ram[3764]  = 1;
  ram[3765]  = 1;
  ram[3766]  = 1;
  ram[3767]  = 1;
  ram[3768]  = 1;
  ram[3769]  = 1;
  ram[3770]  = 1;
  ram[3771]  = 1;
  ram[3772]  = 1;
  ram[3773]  = 1;
  ram[3774]  = 1;
  ram[3775]  = 1;
  ram[3776]  = 1;
  ram[3777]  = 1;
  ram[3778]  = 1;
  ram[3779]  = 1;
  ram[3780]  = 1;
  ram[3781]  = 1;
  ram[3782]  = 1;
  ram[3783]  = 1;
  ram[3784]  = 1;
  ram[3785]  = 1;
  ram[3786]  = 1;
  ram[3787]  = 1;
  ram[3788]  = 1;
  ram[3789]  = 1;
  ram[3790]  = 1;
  ram[3791]  = 1;
  ram[3792]  = 1;
  ram[3793]  = 1;
  ram[3794]  = 1;
  ram[3795]  = 1;
  ram[3796]  = 1;
  ram[3797]  = 1;
  ram[3798]  = 1;
  ram[3799]  = 1;
  ram[3800]  = 1;
  ram[3801]  = 1;
  ram[3802]  = 1;
  ram[3803]  = 1;
  ram[3804]  = 1;
  ram[3805]  = 1;
  ram[3806]  = 1;
  ram[3807]  = 1;
  ram[3808]  = 1;
  ram[3809]  = 1;
  ram[3810]  = 1;
  ram[3811]  = 1;
  ram[3812]  = 1;
  ram[3813]  = 1;
  ram[3814]  = 1;
  ram[3815]  = 1;
  ram[3816]  = 1;
  ram[3817]  = 1;
  ram[3818]  = 1;
  ram[3819]  = 1;
  ram[3820]  = 1;
  ram[3821]  = 1;
  ram[3822]  = 1;
  ram[3823]  = 1;
  ram[3824]  = 1;
  ram[3825]  = 1;
  ram[3826]  = 1;
  ram[3827]  = 1;
  ram[3828]  = 1;
  ram[3829]  = 1;
  ram[3830]  = 1;
  ram[3831]  = 1;
  ram[3832]  = 1;
  ram[3833]  = 1;
  ram[3834]  = 1;
  ram[3835]  = 1;
  ram[3836]  = 1;
  ram[3837]  = 1;
  ram[3838]  = 1;
  ram[3839]  = 1;
  ram[3840]  = 1;
  ram[3841]  = 1;
  ram[3842]  = 1;
  ram[3843]  = 1;
  ram[3844]  = 1;
  ram[3845]  = 1;
  ram[3846]  = 1;
  ram[3847]  = 1;
  ram[3848]  = 1;
  ram[3849]  = 1;
  ram[3850]  = 1;
  ram[3851]  = 1;
  ram[3852]  = 1;
  ram[3853]  = 1;
  ram[3854]  = 1;
  ram[3855]  = 1;
  ram[3856]  = 1;
  ram[3857]  = 1;
  ram[3858]  = 1;
  ram[3859]  = 1;
  ram[3860]  = 1;
  ram[3861]  = 1;
  ram[3862]  = 1;
  ram[3863]  = 1;
  ram[3864]  = 1;
  ram[3865]  = 1;
  ram[3866]  = 1;
  ram[3867]  = 1;
  ram[3868]  = 1;
  ram[3869]  = 1;
  ram[3870]  = 1;
  ram[3871]  = 1;
  ram[3872]  = 1;
  ram[3873]  = 1;
  ram[3874]  = 1;
  ram[3875]  = 1;
  ram[3876]  = 1;
  ram[3877]  = 1;
  ram[3878]  = 1;
  ram[3879]  = 1;
  ram[3880]  = 1;
  ram[3881]  = 1;
  ram[3882]  = 1;
  ram[3883]  = 1;
  ram[3884]  = 1;
  ram[3885]  = 1;
  ram[3886]  = 1;
  ram[3887]  = 1;
  ram[3888]  = 1;
  ram[3889]  = 1;
  ram[3890]  = 1;
  ram[3891]  = 1;
  ram[3892]  = 1;
  ram[3893]  = 1;
  ram[3894]  = 1;
  ram[3895]  = 1;
  ram[3896]  = 1;
  ram[3897]  = 1;
  ram[3898]  = 1;
  ram[3899]  = 1;
  ram[3900]  = 1;
  ram[3901]  = 1;
  ram[3902]  = 1;
  ram[3903]  = 1;
  ram[3904]  = 1;
  ram[3905]  = 1;
  ram[3906]  = 1;
  ram[3907]  = 1;
  ram[3908]  = 1;
  ram[3909]  = 1;
  ram[3910]  = 1;
  ram[3911]  = 1;
  ram[3912]  = 1;
  ram[3913]  = 1;
  ram[3914]  = 1;
  ram[3915]  = 1;
  ram[3916]  = 1;
  ram[3917]  = 1;
  ram[3918]  = 1;
  ram[3919]  = 1;
  ram[3920]  = 1;
  ram[3921]  = 1;
  ram[3922]  = 1;
  ram[3923]  = 1;
  ram[3924]  = 1;
  ram[3925]  = 1;
  ram[3926]  = 1;
  ram[3927]  = 1;
  ram[3928]  = 1;
  ram[3929]  = 1;
  ram[3930]  = 1;
  ram[3931]  = 1;
  ram[3932]  = 1;
  ram[3933]  = 1;
  ram[3934]  = 1;
  ram[3935]  = 1;
  ram[3936]  = 1;
  ram[3937]  = 1;
  ram[3938]  = 1;
  ram[3939]  = 1;
  ram[3940]  = 1;
  ram[3941]  = 1;
  ram[3942]  = 1;
  ram[3943]  = 1;
  ram[3944]  = 1;
  ram[3945]  = 1;
  ram[3946]  = 1;
  ram[3947]  = 1;
  ram[3948]  = 1;
  ram[3949]  = 1;
  ram[3950]  = 1;
  ram[3951]  = 1;
  ram[3952]  = 1;
  ram[3953]  = 1;
  ram[3954]  = 1;
  ram[3955]  = 1;
  ram[3956]  = 1;
  ram[3957]  = 1;
  ram[3958]  = 1;
  ram[3959]  = 1;
  ram[3960]  = 1;
  ram[3961]  = 1;
  ram[3962]  = 1;
  ram[3963]  = 1;
  ram[3964]  = 1;
  ram[3965]  = 1;
  ram[3966]  = 1;
  ram[3967]  = 1;
  ram[3968]  = 1;
  ram[3969]  = 1;
  ram[3970]  = 1;
  ram[3971]  = 1;
  ram[3972]  = 1;
  ram[3973]  = 1;
  ram[3974]  = 1;
  ram[3975]  = 1;
  ram[3976]  = 1;
  ram[3977]  = 1;
  ram[3978]  = 1;
  ram[3979]  = 1;
  ram[3980]  = 1;
  ram[3981]  = 1;
  ram[3982]  = 1;
  ram[3983]  = 1;
  ram[3984]  = 1;
  ram[3985]  = 1;
  ram[3986]  = 1;
  ram[3987]  = 1;
  ram[3988]  = 1;
  ram[3989]  = 1;
  ram[3990]  = 1;
  ram[3991]  = 1;
  ram[3992]  = 1;
  ram[3993]  = 1;
  ram[3994]  = 1;
  ram[3995]  = 1;
  ram[3996]  = 1;
  ram[3997]  = 1;
  ram[3998]  = 1;
  ram[3999]  = 1;
  ram[4000]  = 1;
  ram[4001]  = 1;
  ram[4002]  = 1;
  ram[4003]  = 1;
  ram[4004]  = 1;
  ram[4005]  = 1;
  ram[4006]  = 1;
  ram[4007]  = 1;
  ram[4008]  = 1;
  ram[4009]  = 1;
  ram[4010]  = 1;
  ram[4011]  = 1;
  ram[4012]  = 1;
  ram[4013]  = 1;
  ram[4014]  = 1;
  ram[4015]  = 1;
  ram[4016]  = 1;
  ram[4017]  = 1;
  ram[4018]  = 1;
  ram[4019]  = 1;
  ram[4020]  = 1;
  ram[4021]  = 1;
  ram[4022]  = 1;
  ram[4023]  = 1;
  ram[4024]  = 1;
  ram[4025]  = 1;
  ram[4026]  = 1;
  ram[4027]  = 1;
  ram[4028]  = 1;
  ram[4029]  = 1;
  ram[4030]  = 1;
  ram[4031]  = 1;
  ram[4032]  = 1;
  ram[4033]  = 1;
  ram[4034]  = 1;
  ram[4035]  = 1;
  ram[4036]  = 1;
  ram[4037]  = 1;
  ram[4038]  = 1;
  ram[4039]  = 1;
  ram[4040]  = 1;
  ram[4041]  = 1;
  ram[4042]  = 1;
  ram[4043]  = 1;
  ram[4044]  = 1;
  ram[4045]  = 1;
  ram[4046]  = 1;
  ram[4047]  = 1;
  ram[4048]  = 1;
  ram[4049]  = 1;
  ram[4050]  = 1;
  ram[4051]  = 1;
  ram[4052]  = 1;
  ram[4053]  = 1;
  ram[4054]  = 1;
  ram[4055]  = 1;
  ram[4056]  = 1;
  ram[4057]  = 1;
  ram[4058]  = 1;
  ram[4059]  = 1;
  ram[4060]  = 1;
  ram[4061]  = 1;
  ram[4062]  = 1;
  ram[4063]  = 1;
  ram[4064]  = 1;
  ram[4065]  = 1;
  ram[4066]  = 1;
  ram[4067]  = 1;
  ram[4068]  = 1;
  ram[4069]  = 1;
  ram[4070]  = 1;
  ram[4071]  = 1;
  ram[4072]  = 1;
  ram[4073]  = 1;
  ram[4074]  = 1;
  ram[4075]  = 1;
  ram[4076]  = 1;
  ram[4077]  = 1;
  ram[4078]  = 1;
  ram[4079]  = 1;
  ram[4080]  = 1;
  ram[4081]  = 1;
  ram[4082]  = 1;
  ram[4083]  = 1;
  ram[4084]  = 1;
  ram[4085]  = 1;
  ram[4086]  = 1;
  ram[4087]  = 1;
  ram[4088]  = 1;
  ram[4089]  = 1;
  ram[4090]  = 1;
  ram[4091]  = 1;
  ram[4092]  = 1;
  ram[4093]  = 1;
  ram[4094]  = 1;
  ram[4095]  = 1;
  ram[4096]  = 1;
  ram[4097]  = 1;
  ram[4098]  = 1;
  ram[4099]  = 1;
  ram[4100]  = 1;
  ram[4101]  = 1;
  ram[4102]  = 1;
  ram[4103]  = 1;
  ram[4104]  = 1;
  ram[4105]  = 1;
  ram[4106]  = 1;
  ram[4107]  = 1;
  ram[4108]  = 1;
  ram[4109]  = 1;
  ram[4110]  = 1;
  ram[4111]  = 1;
  ram[4112]  = 1;
  ram[4113]  = 1;
  ram[4114]  = 1;
  ram[4115]  = 1;
  ram[4116]  = 1;
  ram[4117]  = 1;
  ram[4118]  = 1;
  ram[4119]  = 1;
  ram[4120]  = 1;
  ram[4121]  = 1;
  ram[4122]  = 1;
  ram[4123]  = 1;
  ram[4124]  = 1;
  ram[4125]  = 1;
  ram[4126]  = 1;
  ram[4127]  = 1;
  ram[4128]  = 1;
  ram[4129]  = 1;
  ram[4130]  = 1;
  ram[4131]  = 1;
  ram[4132]  = 1;
  ram[4133]  = 1;
  ram[4134]  = 1;
  ram[4135]  = 1;
  ram[4136]  = 1;
  ram[4137]  = 1;
  ram[4138]  = 1;
  ram[4139]  = 1;
  ram[4140]  = 1;
  ram[4141]  = 1;
  ram[4142]  = 1;
  ram[4143]  = 1;
  ram[4144]  = 1;
  ram[4145]  = 1;
  ram[4146]  = 1;
  ram[4147]  = 1;
  ram[4148]  = 1;
  ram[4149]  = 1;
  ram[4150]  = 1;
  ram[4151]  = 1;
  ram[4152]  = 1;
  ram[4153]  = 1;
  ram[4154]  = 1;
  ram[4155]  = 1;
  ram[4156]  = 1;
  ram[4157]  = 1;
  ram[4158]  = 1;
  ram[4159]  = 1;
  ram[4160]  = 1;
  ram[4161]  = 1;
  ram[4162]  = 1;
  ram[4163]  = 1;
  ram[4164]  = 1;
  ram[4165]  = 1;
  ram[4166]  = 1;
  ram[4167]  = 1;
  ram[4168]  = 1;
  ram[4169]  = 1;
  ram[4170]  = 1;
  ram[4171]  = 1;
  ram[4172]  = 1;
  ram[4173]  = 1;
  ram[4174]  = 1;
  ram[4175]  = 1;
  ram[4176]  = 1;
  ram[4177]  = 1;
  ram[4178]  = 1;
  ram[4179]  = 1;
  ram[4180]  = 1;
  ram[4181]  = 1;
  ram[4182]  = 1;
  ram[4183]  = 1;
  ram[4184]  = 1;
  ram[4185]  = 1;
  ram[4186]  = 1;
  ram[4187]  = 1;
  ram[4188]  = 1;
  ram[4189]  = 1;
  ram[4190]  = 1;
  ram[4191]  = 1;
  ram[4192]  = 1;
  ram[4193]  = 1;
  ram[4194]  = 1;
  ram[4195]  = 1;
  ram[4196]  = 1;
  ram[4197]  = 1;
  ram[4198]  = 1;
  ram[4199]  = 1;
  ram[4200]  = 1;
  ram[4201]  = 1;
  ram[4202]  = 1;
  ram[4203]  = 1;
  ram[4204]  = 1;
  ram[4205]  = 1;
  ram[4206]  = 1;
  ram[4207]  = 1;
  ram[4208]  = 1;
  ram[4209]  = 1;
  ram[4210]  = 1;
  ram[4211]  = 1;
  ram[4212]  = 1;
  ram[4213]  = 1;
  ram[4214]  = 1;
  ram[4215]  = 1;
  ram[4216]  = 1;
  ram[4217]  = 1;
  ram[4218]  = 1;
  ram[4219]  = 1;
  ram[4220]  = 1;
  ram[4221]  = 1;
  ram[4222]  = 1;
  ram[4223]  = 1;
  ram[4224]  = 1;
  ram[4225]  = 1;
  ram[4226]  = 1;
  ram[4227]  = 1;
  ram[4228]  = 1;
  ram[4229]  = 1;
  ram[4230]  = 1;
  ram[4231]  = 1;
  ram[4232]  = 1;
  ram[4233]  = 1;
  ram[4234]  = 1;
  ram[4235]  = 1;
  ram[4236]  = 1;
  ram[4237]  = 1;
  ram[4238]  = 1;
  ram[4239]  = 1;
  ram[4240]  = 1;
  ram[4241]  = 1;
  ram[4242]  = 1;
  ram[4243]  = 1;
  ram[4244]  = 1;
  ram[4245]  = 1;
  ram[4246]  = 1;
  ram[4247]  = 1;
  ram[4248]  = 1;
  ram[4249]  = 1;
  ram[4250]  = 1;
  ram[4251]  = 1;
  ram[4252]  = 1;
  ram[4253]  = 1;
  ram[4254]  = 1;
  ram[4255]  = 1;
  ram[4256]  = 1;
  ram[4257]  = 1;
  ram[4258]  = 1;
  ram[4259]  = 1;
  ram[4260]  = 1;
  ram[4261]  = 1;
  ram[4262]  = 1;
  ram[4263]  = 1;
  ram[4264]  = 1;
  ram[4265]  = 1;
  ram[4266]  = 1;
  ram[4267]  = 1;
  ram[4268]  = 1;
  ram[4269]  = 1;
  ram[4270]  = 1;
  ram[4271]  = 1;
  ram[4272]  = 1;
  ram[4273]  = 1;
  ram[4274]  = 1;
  ram[4275]  = 1;
  ram[4276]  = 1;
  ram[4277]  = 1;
  ram[4278]  = 1;
  ram[4279]  = 1;
  ram[4280]  = 1;
  ram[4281]  = 1;
  ram[4282]  = 1;
  ram[4283]  = 1;
  ram[4284]  = 1;
  ram[4285]  = 1;
  ram[4286]  = 1;
  ram[4287]  = 1;
  ram[4288]  = 1;
  ram[4289]  = 1;
  ram[4290]  = 1;
  ram[4291]  = 1;
  ram[4292]  = 1;
  ram[4293]  = 1;
  ram[4294]  = 1;
  ram[4295]  = 1;
  ram[4296]  = 1;
  ram[4297]  = 1;
  ram[4298]  = 1;
  ram[4299]  = 1;
  ram[4300]  = 1;
  ram[4301]  = 1;
  ram[4302]  = 1;
  ram[4303]  = 1;
  ram[4304]  = 1;
  ram[4305]  = 1;
  ram[4306]  = 1;
  ram[4307]  = 1;
  ram[4308]  = 1;
  ram[4309]  = 1;
  ram[4310]  = 1;
  ram[4311]  = 1;
  ram[4312]  = 1;
  ram[4313]  = 1;
  ram[4314]  = 1;
  ram[4315]  = 1;
  ram[4316]  = 1;
  ram[4317]  = 1;
  ram[4318]  = 1;
  ram[4319]  = 1;
  ram[4320]  = 1;
  ram[4321]  = 1;
  ram[4322]  = 1;
  ram[4323]  = 1;
  ram[4324]  = 1;
  ram[4325]  = 1;
  ram[4326]  = 1;
  ram[4327]  = 1;
  ram[4328]  = 1;
  ram[4329]  = 1;
  ram[4330]  = 1;
  ram[4331]  = 1;
  ram[4332]  = 1;
  ram[4333]  = 1;
  ram[4334]  = 1;
  ram[4335]  = 1;
  ram[4336]  = 1;
  ram[4337]  = 1;
  ram[4338]  = 1;
  ram[4339]  = 1;
  ram[4340]  = 1;
  ram[4341]  = 1;
  ram[4342]  = 1;
  ram[4343]  = 1;
  ram[4344]  = 1;
  ram[4345]  = 1;
  ram[4346]  = 1;
  ram[4347]  = 1;
  ram[4348]  = 1;
  ram[4349]  = 1;
  ram[4350]  = 1;
  ram[4351]  = 1;
  ram[4352]  = 1;
  ram[4353]  = 1;
  ram[4354]  = 1;
  ram[4355]  = 1;
  ram[4356]  = 1;
  ram[4357]  = 1;
  ram[4358]  = 1;
  ram[4359]  = 1;
  ram[4360]  = 1;
  ram[4361]  = 1;
  ram[4362]  = 1;
  ram[4363]  = 1;
  ram[4364]  = 1;
  ram[4365]  = 1;
  ram[4366]  = 1;
  ram[4367]  = 1;
  ram[4368]  = 1;
  ram[4369]  = 1;
  ram[4370]  = 1;
  ram[4371]  = 1;
  ram[4372]  = 1;
  ram[4373]  = 1;
  ram[4374]  = 1;
  ram[4375]  = 1;
  ram[4376]  = 1;
  ram[4377]  = 1;
  ram[4378]  = 1;
  ram[4379]  = 1;
  ram[4380]  = 1;
  ram[4381]  = 1;
  ram[4382]  = 1;
  ram[4383]  = 1;
  ram[4384]  = 1;
  ram[4385]  = 1;
  ram[4386]  = 1;
  ram[4387]  = 1;
  ram[4388]  = 1;
  ram[4389]  = 1;
  ram[4390]  = 1;
  ram[4391]  = 1;
  ram[4392]  = 1;
  ram[4393]  = 1;
  ram[4394]  = 1;
  ram[4395]  = 1;
  ram[4396]  = 1;
  ram[4397]  = 1;
  ram[4398]  = 1;
  ram[4399]  = 1;
  ram[4400]  = 1;
  ram[4401]  = 1;
  ram[4402]  = 1;
  ram[4403]  = 1;
  ram[4404]  = 1;
  ram[4405]  = 1;
  ram[4406]  = 1;
  ram[4407]  = 1;
  ram[4408]  = 1;
  ram[4409]  = 1;
  ram[4410]  = 1;
  ram[4411]  = 1;
  ram[4412]  = 1;
  ram[4413]  = 1;
  ram[4414]  = 1;
  ram[4415]  = 1;
  ram[4416]  = 1;
  ram[4417]  = 1;
  ram[4418]  = 1;
  ram[4419]  = 1;
  ram[4420]  = 1;
  ram[4421]  = 1;
  ram[4422]  = 1;
  ram[4423]  = 1;
  ram[4424]  = 1;
  ram[4425]  = 1;
  ram[4426]  = 1;
  ram[4427]  = 1;
  ram[4428]  = 1;
  ram[4429]  = 1;
  ram[4430]  = 1;
  ram[4431]  = 1;
  ram[4432]  = 1;
  ram[4433]  = 1;
  ram[4434]  = 1;
  ram[4435]  = 1;
  ram[4436]  = 1;
  ram[4437]  = 1;
  ram[4438]  = 1;
  ram[4439]  = 1;
  ram[4440]  = 1;
  ram[4441]  = 1;
  ram[4442]  = 1;
  ram[4443]  = 1;
  ram[4444]  = 1;
  ram[4445]  = 1;
  ram[4446]  = 1;
  ram[4447]  = 1;
  ram[4448]  = 1;
  ram[4449]  = 1;
  ram[4450]  = 1;
  ram[4451]  = 1;
  ram[4452]  = 1;
  ram[4453]  = 1;
  ram[4454]  = 1;
  ram[4455]  = 1;
  ram[4456]  = 1;
  ram[4457]  = 1;
  ram[4458]  = 1;
  ram[4459]  = 1;
  ram[4460]  = 1;
  ram[4461]  = 1;
  ram[4462]  = 1;
  ram[4463]  = 1;
  ram[4464]  = 1;
  ram[4465]  = 1;
  ram[4466]  = 1;
  ram[4467]  = 1;
  ram[4468]  = 1;
  ram[4469]  = 1;
  ram[4470]  = 1;
  ram[4471]  = 1;
  ram[4472]  = 1;
  ram[4473]  = 1;
  ram[4474]  = 1;
  ram[4475]  = 1;
  ram[4476]  = 1;
  ram[4477]  = 1;
  ram[4478]  = 1;
  ram[4479]  = 1;
  ram[4480]  = 1;
  ram[4481]  = 1;
  ram[4482]  = 1;
  ram[4483]  = 1;
  ram[4484]  = 1;
  ram[4485]  = 1;
  ram[4486]  = 1;
  ram[4487]  = 1;
  ram[4488]  = 1;
  ram[4489]  = 1;
  ram[4490]  = 1;
  ram[4491]  = 1;
  ram[4492]  = 1;
  ram[4493]  = 1;
  ram[4494]  = 1;
  ram[4495]  = 1;
  ram[4496]  = 1;
  ram[4497]  = 1;
  ram[4498]  = 1;
  ram[4499]  = 1;
  ram[4500]  = 1;
  ram[4501]  = 1;
  ram[4502]  = 1;
  ram[4503]  = 1;
  ram[4504]  = 1;
  ram[4505]  = 1;
  ram[4506]  = 1;
  ram[4507]  = 1;
  ram[4508]  = 1;
  ram[4509]  = 1;
  ram[4510]  = 1;
  ram[4511]  = 1;
  ram[4512]  = 1;
  ram[4513]  = 1;
  ram[4514]  = 1;
  ram[4515]  = 1;
  ram[4516]  = 1;
  ram[4517]  = 1;
  ram[4518]  = 1;
  ram[4519]  = 1;
  ram[4520]  = 1;
  ram[4521]  = 1;
  ram[4522]  = 1;
  ram[4523]  = 1;
  ram[4524]  = 1;
  ram[4525]  = 1;
  ram[4526]  = 1;
  ram[4527]  = 1;
  ram[4528]  = 1;
  ram[4529]  = 1;
  ram[4530]  = 1;
  ram[4531]  = 1;
  ram[4532]  = 1;
  ram[4533]  = 1;
  ram[4534]  = 1;
  ram[4535]  = 1;
  ram[4536]  = 1;
  ram[4537]  = 1;
  ram[4538]  = 1;
  ram[4539]  = 1;
  ram[4540]  = 1;
  ram[4541]  = 1;
  ram[4542]  = 1;
  ram[4543]  = 1;
  ram[4544]  = 1;
  ram[4545]  = 1;
  ram[4546]  = 1;
  ram[4547]  = 1;
  ram[4548]  = 1;
  ram[4549]  = 1;
  ram[4550]  = 1;
  ram[4551]  = 1;
  ram[4552]  = 1;
  ram[4553]  = 1;
  ram[4554]  = 1;
  ram[4555]  = 1;
  ram[4556]  = 1;
  ram[4557]  = 1;
  ram[4558]  = 1;
  ram[4559]  = 1;
  ram[4560]  = 1;
  ram[4561]  = 1;
  ram[4562]  = 1;
  ram[4563]  = 1;
  ram[4564]  = 1;
  ram[4565]  = 1;
  ram[4566]  = 1;
  ram[4567]  = 1;
  ram[4568]  = 1;
  ram[4569]  = 1;
  ram[4570]  = 1;
  ram[4571]  = 1;
  ram[4572]  = 1;
  ram[4573]  = 1;
  ram[4574]  = 1;
  ram[4575]  = 1;
  ram[4576]  = 1;
  ram[4577]  = 1;
  ram[4578]  = 1;
  ram[4579]  = 1;
  ram[4580]  = 1;
  ram[4581]  = 1;
  ram[4582]  = 1;
  ram[4583]  = 1;
  ram[4584]  = 1;
  ram[4585]  = 1;
  ram[4586]  = 1;
  ram[4587]  = 1;
  ram[4588]  = 1;
  ram[4589]  = 1;
  ram[4590]  = 1;
  ram[4591]  = 1;
  ram[4592]  = 1;
  ram[4593]  = 1;
  ram[4594]  = 1;
  ram[4595]  = 1;
  ram[4596]  = 1;
  ram[4597]  = 1;
  ram[4598]  = 1;
  ram[4599]  = 1;
  ram[4600]  = 1;
  ram[4601]  = 1;
  ram[4602]  = 1;
  ram[4603]  = 1;
  ram[4604]  = 1;
  ram[4605]  = 1;
  ram[4606]  = 1;
  ram[4607]  = 1;
  ram[4608]  = 1;
  ram[4609]  = 1;
  ram[4610]  = 1;
  ram[4611]  = 1;
  ram[4612]  = 1;
  ram[4613]  = 1;
  ram[4614]  = 1;
  ram[4615]  = 1;
  ram[4616]  = 1;
  ram[4617]  = 1;
  ram[4618]  = 1;
  ram[4619]  = 1;
  ram[4620]  = 1;
  ram[4621]  = 1;
  ram[4622]  = 1;
  ram[4623]  = 1;
  ram[4624]  = 1;
  ram[4625]  = 1;
  ram[4626]  = 1;
  ram[4627]  = 1;
  ram[4628]  = 1;
  ram[4629]  = 1;
  ram[4630]  = 1;
  ram[4631]  = 1;
  ram[4632]  = 1;
  ram[4633]  = 1;
  ram[4634]  = 1;
  ram[4635]  = 1;
  ram[4636]  = 1;
  ram[4637]  = 1;
  ram[4638]  = 1;
  ram[4639]  = 1;
  ram[4640]  = 1;
  ram[4641]  = 1;
  ram[4642]  = 1;
  ram[4643]  = 1;
  ram[4644]  = 1;
  ram[4645]  = 1;
  ram[4646]  = 1;
  ram[4647]  = 1;
  ram[4648]  = 1;
  ram[4649]  = 1;
  ram[4650]  = 1;
  ram[4651]  = 1;
  ram[4652]  = 1;
  ram[4653]  = 1;
  ram[4654]  = 1;
  ram[4655]  = 1;
  ram[4656]  = 1;
  ram[4657]  = 1;
  ram[4658]  = 1;
  ram[4659]  = 1;
  ram[4660]  = 1;
  ram[4661]  = 1;
  ram[4662]  = 1;
  ram[4663]  = 1;
  ram[4664]  = 1;
  ram[4665]  = 1;
  ram[4666]  = 1;
  ram[4667]  = 1;
  ram[4668]  = 1;
  ram[4669]  = 1;
  ram[4670]  = 1;
  ram[4671]  = 1;
  ram[4672]  = 1;
  ram[4673]  = 1;
  ram[4674]  = 1;
  ram[4675]  = 1;
  ram[4676]  = 1;
  ram[4677]  = 1;
  ram[4678]  = 1;
  ram[4679]  = 1;
  ram[4680]  = 1;
  ram[4681]  = 1;
  ram[4682]  = 1;
  ram[4683]  = 1;
  ram[4684]  = 1;
  ram[4685]  = 1;
  ram[4686]  = 1;
  ram[4687]  = 1;
  ram[4688]  = 1;
  ram[4689]  = 1;
  ram[4690]  = 1;
  ram[4691]  = 1;
  ram[4692]  = 1;
  ram[4693]  = 1;
  ram[4694]  = 1;
  ram[4695]  = 1;
  ram[4696]  = 1;
  ram[4697]  = 1;
  ram[4698]  = 1;
  ram[4699]  = 1;
  ram[4700]  = 1;
  ram[4701]  = 1;
  ram[4702]  = 1;
  ram[4703]  = 1;
  ram[4704]  = 1;
  ram[4705]  = 1;
  ram[4706]  = 1;
  ram[4707]  = 1;
  ram[4708]  = 1;
  ram[4709]  = 1;
  ram[4710]  = 1;
  ram[4711]  = 1;
  ram[4712]  = 1;
  ram[4713]  = 1;
  ram[4714]  = 1;
  ram[4715]  = 1;
  ram[4716]  = 1;
  ram[4717]  = 1;
  ram[4718]  = 1;
  ram[4719]  = 1;
  ram[4720]  = 1;
  ram[4721]  = 1;
  ram[4722]  = 1;
  ram[4723]  = 1;
  ram[4724]  = 1;
  ram[4725]  = 1;
  ram[4726]  = 1;
  ram[4727]  = 1;
  ram[4728]  = 1;
  ram[4729]  = 1;
  ram[4730]  = 1;
  ram[4731]  = 1;
  ram[4732]  = 1;
  ram[4733]  = 1;
  ram[4734]  = 1;
  ram[4735]  = 1;
  ram[4736]  = 1;
  ram[4737]  = 1;
  ram[4738]  = 1;
  ram[4739]  = 1;
  ram[4740]  = 1;
  ram[4741]  = 1;
  ram[4742]  = 1;
  ram[4743]  = 1;
  ram[4744]  = 1;
  ram[4745]  = 1;
  ram[4746]  = 1;
  ram[4747]  = 1;
  ram[4748]  = 1;
  ram[4749]  = 1;
  ram[4750]  = 1;
  ram[4751]  = 1;
  ram[4752]  = 1;
  ram[4753]  = 1;
  ram[4754]  = 1;
  ram[4755]  = 1;
  ram[4756]  = 1;
  ram[4757]  = 1;
  ram[4758]  = 1;
  ram[4759]  = 1;
  ram[4760]  = 1;
  ram[4761]  = 1;
  ram[4762]  = 1;
  ram[4763]  = 1;
  ram[4764]  = 1;
  ram[4765]  = 1;
  ram[4766]  = 1;
  ram[4767]  = 1;
  ram[4768]  = 1;
  ram[4769]  = 1;
  ram[4770]  = 1;
  ram[4771]  = 1;
  ram[4772]  = 1;
  ram[4773]  = 1;
  ram[4774]  = 1;
  ram[4775]  = 1;
  ram[4776]  = 1;
  ram[4777]  = 1;
  ram[4778]  = 1;
  ram[4779]  = 1;
  ram[4780]  = 1;
  ram[4781]  = 1;
  ram[4782]  = 1;
  ram[4783]  = 1;
  ram[4784]  = 1;
  ram[4785]  = 1;
  ram[4786]  = 1;
  ram[4787]  = 1;
  ram[4788]  = 1;
  ram[4789]  = 1;
  ram[4790]  = 1;
  ram[4791]  = 1;
  ram[4792]  = 1;
  ram[4793]  = 1;
  ram[4794]  = 1;
  ram[4795]  = 1;
  ram[4796]  = 1;
  ram[4797]  = 1;
  ram[4798]  = 1;
  ram[4799]  = 1;
  ram[4800]  = 1;
  ram[4801]  = 1;
  ram[4802]  = 1;
  ram[4803]  = 1;
  ram[4804]  = 1;
  ram[4805]  = 1;
  ram[4806]  = 1;
  ram[4807]  = 1;
  ram[4808]  = 1;
  ram[4809]  = 1;
  ram[4810]  = 1;
  ram[4811]  = 1;
  ram[4812]  = 1;
  ram[4813]  = 1;
  ram[4814]  = 1;
  ram[4815]  = 1;
  ram[4816]  = 1;
  ram[4817]  = 1;
  ram[4818]  = 1;
  ram[4819]  = 1;
  ram[4820]  = 1;
  ram[4821]  = 1;
  ram[4822]  = 1;
  ram[4823]  = 1;
  ram[4824]  = 1;
  ram[4825]  = 1;
  ram[4826]  = 1;
  ram[4827]  = 1;
  ram[4828]  = 1;
  ram[4829]  = 1;
  ram[4830]  = 1;
  ram[4831]  = 1;
  ram[4832]  = 1;
  ram[4833]  = 1;
  ram[4834]  = 1;
  ram[4835]  = 1;
  ram[4836]  = 1;
  ram[4837]  = 1;
  ram[4838]  = 1;
  ram[4839]  = 1;
  ram[4840]  = 1;
  ram[4841]  = 1;
  ram[4842]  = 1;
  ram[4843]  = 1;
  ram[4844]  = 1;
  ram[4845]  = 1;
  ram[4846]  = 1;
  ram[4847]  = 1;
  ram[4848]  = 1;
  ram[4849]  = 1;
  ram[4850]  = 1;
  ram[4851]  = 1;
  ram[4852]  = 1;
  ram[4853]  = 1;
  ram[4854]  = 1;
  ram[4855]  = 1;
  ram[4856]  = 1;
  ram[4857]  = 1;
  ram[4858]  = 1;
  ram[4859]  = 1;
  ram[4860]  = 1;
  ram[4861]  = 1;
  ram[4862]  = 1;
  ram[4863]  = 1;
  ram[4864]  = 1;
  ram[4865]  = 1;
  ram[4866]  = 1;
  ram[4867]  = 1;
  ram[4868]  = 1;
  ram[4869]  = 1;
  ram[4870]  = 1;
  ram[4871]  = 1;
  ram[4872]  = 1;
  ram[4873]  = 1;
  ram[4874]  = 1;
  ram[4875]  = 1;
  ram[4876]  = 1;
  ram[4877]  = 1;
  ram[4878]  = 1;
  ram[4879]  = 1;
  ram[4880]  = 1;
  ram[4881]  = 1;
  ram[4882]  = 1;
  ram[4883]  = 1;
  ram[4884]  = 1;
  ram[4885]  = 1;
  ram[4886]  = 1;
  ram[4887]  = 1;
  ram[4888]  = 1;
  ram[4889]  = 1;
  ram[4890]  = 1;
  ram[4891]  = 1;
  ram[4892]  = 1;
  ram[4893]  = 1;
  ram[4894]  = 1;
  ram[4895]  = 1;
  ram[4896]  = 1;
  ram[4897]  = 1;
  ram[4898]  = 1;
  ram[4899]  = 1;
  ram[4900]  = 1;
  ram[4901]  = 1;
  ram[4902]  = 1;
  ram[4903]  = 1;
  ram[4904]  = 1;
  ram[4905]  = 1;
  ram[4906]  = 1;
  ram[4907]  = 1;
  ram[4908]  = 1;
  ram[4909]  = 1;
  ram[4910]  = 1;
  ram[4911]  = 1;
  ram[4912]  = 1;
  ram[4913]  = 1;
  ram[4914]  = 1;
  ram[4915]  = 1;
  ram[4916]  = 1;
  ram[4917]  = 1;
  ram[4918]  = 1;
  ram[4919]  = 1;
  ram[4920]  = 1;
  ram[4921]  = 1;
  ram[4922]  = 1;
  ram[4923]  = 1;
  ram[4924]  = 1;
  ram[4925]  = 1;
  ram[4926]  = 1;
  ram[4927]  = 1;
  ram[4928]  = 1;
  ram[4929]  = 1;
  ram[4930]  = 1;
  ram[4931]  = 1;
  ram[4932]  = 1;
  ram[4933]  = 1;
  ram[4934]  = 1;
  ram[4935]  = 1;
  ram[4936]  = 1;
  ram[4937]  = 1;
  ram[4938]  = 1;
  ram[4939]  = 1;
  ram[4940]  = 1;
  ram[4941]  = 1;
  ram[4942]  = 1;
  ram[4943]  = 1;
  ram[4944]  = 1;
  ram[4945]  = 1;
  ram[4946]  = 1;
  ram[4947]  = 1;
  ram[4948]  = 1;
  ram[4949]  = 1;
  ram[4950]  = 1;
  ram[4951]  = 1;
  ram[4952]  = 1;
  ram[4953]  = 1;
  ram[4954]  = 1;
  ram[4955]  = 1;
  ram[4956]  = 1;
  ram[4957]  = 1;
  ram[4958]  = 1;
  ram[4959]  = 1;
  ram[4960]  = 1;
  ram[4961]  = 1;
  ram[4962]  = 1;
  ram[4963]  = 1;
  ram[4964]  = 1;
  ram[4965]  = 1;
  ram[4966]  = 1;
  ram[4967]  = 1;
  ram[4968]  = 1;
  ram[4969]  = 1;
  ram[4970]  = 1;
  ram[4971]  = 1;
  ram[4972]  = 1;
  ram[4973]  = 1;
  ram[4974]  = 1;
  ram[4975]  = 1;
  ram[4976]  = 1;
  ram[4977]  = 1;
  ram[4978]  = 1;
  ram[4979]  = 1;
  ram[4980]  = 1;
  ram[4981]  = 1;
  ram[4982]  = 1;
  ram[4983]  = 1;
  ram[4984]  = 1;
  ram[4985]  = 1;
  ram[4986]  = 1;
  ram[4987]  = 1;
  ram[4988]  = 1;
  ram[4989]  = 1;
  ram[4990]  = 1;
  ram[4991]  = 1;
  ram[4992]  = 1;
  ram[4993]  = 1;
  ram[4994]  = 1;
  ram[4995]  = 1;
  ram[4996]  = 1;
  ram[4997]  = 1;
  ram[4998]  = 1;
  ram[4999]  = 1;
  ram[5000]  = 1;
  ram[5001]  = 1;
  ram[5002]  = 1;
  ram[5003]  = 1;
  ram[5004]  = 1;
  ram[5005]  = 1;
  ram[5006]  = 1;
  ram[5007]  = 1;
  ram[5008]  = 1;
  ram[5009]  = 1;
  ram[5010]  = 1;
  ram[5011]  = 1;
  ram[5012]  = 1;
  ram[5013]  = 1;
  ram[5014]  = 1;
  ram[5015]  = 1;
  ram[5016]  = 1;
  ram[5017]  = 1;
  ram[5018]  = 1;
  ram[5019]  = 1;
  ram[5020]  = 1;
  ram[5021]  = 1;
  ram[5022]  = 1;
  ram[5023]  = 1;
  ram[5024]  = 1;
  ram[5025]  = 1;
  ram[5026]  = 1;
  ram[5027]  = 1;
  ram[5028]  = 1;
  ram[5029]  = 1;
  ram[5030]  = 1;
  ram[5031]  = 1;
  ram[5032]  = 1;
  ram[5033]  = 1;
  ram[5034]  = 1;
  ram[5035]  = 1;
  ram[5036]  = 1;
  ram[5037]  = 1;
  ram[5038]  = 1;
  ram[5039]  = 1;
  ram[5040]  = 1;
  ram[5041]  = 1;
  ram[5042]  = 1;
  ram[5043]  = 1;
  ram[5044]  = 1;
  ram[5045]  = 1;
  ram[5046]  = 1;
  ram[5047]  = 1;
  ram[5048]  = 1;
  ram[5049]  = 1;
  ram[5050]  = 1;
  ram[5051]  = 1;
  ram[5052]  = 1;
  ram[5053]  = 1;
  ram[5054]  = 1;
  ram[5055]  = 1;
  ram[5056]  = 1;
  ram[5057]  = 1;
  ram[5058]  = 1;
  ram[5059]  = 1;
  ram[5060]  = 1;
  ram[5061]  = 1;
  ram[5062]  = 1;
  ram[5063]  = 1;
  ram[5064]  = 1;
  ram[5065]  = 1;
  ram[5066]  = 1;
  ram[5067]  = 1;
  ram[5068]  = 1;
  ram[5069]  = 1;
  ram[5070]  = 1;
  ram[5071]  = 1;
  ram[5072]  = 1;
  ram[5073]  = 1;
  ram[5074]  = 1;
  ram[5075]  = 1;
  ram[5076]  = 1;
  ram[5077]  = 1;
  ram[5078]  = 1;
  ram[5079]  = 1;
  ram[5080]  = 1;
  ram[5081]  = 1;
  ram[5082]  = 1;
  ram[5083]  = 1;
  ram[5084]  = 1;
  ram[5085]  = 1;
  ram[5086]  = 1;
  ram[5087]  = 1;
  ram[5088]  = 1;
  ram[5089]  = 1;
  ram[5090]  = 1;
  ram[5091]  = 1;
  ram[5092]  = 1;
  ram[5093]  = 1;
  ram[5094]  = 1;
  ram[5095]  = 1;
  ram[5096]  = 1;
  ram[5097]  = 1;
  ram[5098]  = 1;
  ram[5099]  = 1;
  ram[5100]  = 1;
  ram[5101]  = 1;
  ram[5102]  = 1;
  ram[5103]  = 1;
  ram[5104]  = 1;
  ram[5105]  = 1;
  ram[5106]  = 1;
  ram[5107]  = 1;
  ram[5108]  = 1;
  ram[5109]  = 1;
  ram[5110]  = 1;
  ram[5111]  = 1;
  ram[5112]  = 1;
  ram[5113]  = 1;
  ram[5114]  = 1;
  ram[5115]  = 1;
  ram[5116]  = 1;
  ram[5117]  = 1;
  ram[5118]  = 1;
  ram[5119]  = 1;
  ram[5120]  = 1;
  ram[5121]  = 1;
  ram[5122]  = 1;
  ram[5123]  = 1;
  ram[5124]  = 1;
  ram[5125]  = 1;
  ram[5126]  = 1;
  ram[5127]  = 1;
  ram[5128]  = 1;
  ram[5129]  = 1;
  ram[5130]  = 1;
  ram[5131]  = 1;
  ram[5132]  = 1;
  ram[5133]  = 1;
  ram[5134]  = 1;
  ram[5135]  = 1;
  ram[5136]  = 1;
  ram[5137]  = 1;
  ram[5138]  = 1;
  ram[5139]  = 1;
  ram[5140]  = 1;
  ram[5141]  = 1;
  ram[5142]  = 1;
  ram[5143]  = 1;
  ram[5144]  = 1;
  ram[5145]  = 1;
  ram[5146]  = 1;
  ram[5147]  = 1;
  ram[5148]  = 1;
  ram[5149]  = 1;
  ram[5150]  = 1;
  ram[5151]  = 1;
  ram[5152]  = 1;
  ram[5153]  = 1;
  ram[5154]  = 1;
  ram[5155]  = 1;
  ram[5156]  = 1;
  ram[5157]  = 1;
  ram[5158]  = 1;
  ram[5159]  = 1;
  ram[5160]  = 1;
  ram[5161]  = 1;
  ram[5162]  = 1;
  ram[5163]  = 1;
  ram[5164]  = 1;
  ram[5165]  = 1;
  ram[5166]  = 1;
  ram[5167]  = 1;
  ram[5168]  = 1;
  ram[5169]  = 1;
  ram[5170]  = 1;
  ram[5171]  = 1;
  ram[5172]  = 1;
  ram[5173]  = 1;
  ram[5174]  = 1;
  ram[5175]  = 1;
  ram[5176]  = 1;
  ram[5177]  = 1;
  ram[5178]  = 1;
  ram[5179]  = 1;
  ram[5180]  = 1;
  ram[5181]  = 1;
  ram[5182]  = 1;
  ram[5183]  = 1;
  ram[5184]  = 1;
  ram[5185]  = 1;
  ram[5186]  = 1;
  ram[5187]  = 1;
  ram[5188]  = 1;
  ram[5189]  = 1;
  ram[5190]  = 1;
  ram[5191]  = 1;
  ram[5192]  = 1;
  ram[5193]  = 1;
  ram[5194]  = 1;
  ram[5195]  = 1;
  ram[5196]  = 1;
  ram[5197]  = 1;
  ram[5198]  = 1;
  ram[5199]  = 1;
  ram[5200]  = 1;
  ram[5201]  = 1;
  ram[5202]  = 1;
  ram[5203]  = 0;
  ram[5204]  = 0;
  ram[5205]  = 0;
  ram[5206]  = 0;
  ram[5207]  = 0;
  ram[5208]  = 1;
  ram[5209]  = 1;
  ram[5210]  = 1;
  ram[5211]  = 1;
  ram[5212]  = 1;
  ram[5213]  = 1;
  ram[5214]  = 1;
  ram[5215]  = 1;
  ram[5216]  = 1;
  ram[5217]  = 1;
  ram[5218]  = 1;
  ram[5219]  = 1;
  ram[5220]  = 1;
  ram[5221]  = 1;
  ram[5222]  = 1;
  ram[5223]  = 1;
  ram[5224]  = 1;
  ram[5225]  = 1;
  ram[5226]  = 1;
  ram[5227]  = 1;
  ram[5228]  = 1;
  ram[5229]  = 1;
  ram[5230]  = 1;
  ram[5231]  = 1;
  ram[5232]  = 1;
  ram[5233]  = 1;
  ram[5234]  = 1;
  ram[5235]  = 1;
  ram[5236]  = 1;
  ram[5237]  = 1;
  ram[5238]  = 1;
  ram[5239]  = 1;
  ram[5240]  = 1;
  ram[5241]  = 1;
  ram[5242]  = 1;
  ram[5243]  = 1;
  ram[5244]  = 1;
  ram[5245]  = 1;
  ram[5246]  = 1;
  ram[5247]  = 1;
  ram[5248]  = 1;
  ram[5249]  = 1;
  ram[5250]  = 1;
  ram[5251]  = 1;
  ram[5252]  = 1;
  ram[5253]  = 1;
  ram[5254]  = 1;
  ram[5255]  = 0;
  ram[5256]  = 0;
  ram[5257]  = 0;
  ram[5258]  = 0;
  ram[5259]  = 0;
  ram[5260]  = 0;
  ram[5261]  = 1;
  ram[5262]  = 1;
  ram[5263]  = 1;
  ram[5264]  = 1;
  ram[5265]  = 1;
  ram[5266]  = 1;
  ram[5267]  = 1;
  ram[5268]  = 1;
  ram[5269]  = 1;
  ram[5270]  = 1;
  ram[5271]  = 1;
  ram[5272]  = 1;
  ram[5273]  = 1;
  ram[5274]  = 1;
  ram[5275]  = 1;
  ram[5276]  = 1;
  ram[5277]  = 1;
  ram[5278]  = 1;
  ram[5279]  = 1;
  ram[5280]  = 1;
  ram[5281]  = 1;
  ram[5282]  = 1;
  ram[5283]  = 1;
  ram[5284]  = 1;
  ram[5285]  = 1;
  ram[5286]  = 1;
  ram[5287]  = 1;
  ram[5288]  = 1;
  ram[5289]  = 1;
  ram[5290]  = 1;
  ram[5291]  = 0;
  ram[5292]  = 0;
  ram[5293]  = 1;
  ram[5294]  = 1;
  ram[5295]  = 1;
  ram[5296]  = 1;
  ram[5297]  = 1;
  ram[5298]  = 1;
  ram[5299]  = 1;
  ram[5300]  = 1;
  ram[5301]  = 1;
  ram[5302]  = 1;
  ram[5303]  = 1;
  ram[5304]  = 1;
  ram[5305]  = 1;
  ram[5306]  = 1;
  ram[5307]  = 1;
  ram[5308]  = 1;
  ram[5309]  = 1;
  ram[5310]  = 1;
  ram[5311]  = 1;
  ram[5312]  = 1;
  ram[5313]  = 1;
  ram[5314]  = 1;
  ram[5315]  = 1;
  ram[5316]  = 1;
  ram[5317]  = 1;
  ram[5318]  = 1;
  ram[5319]  = 1;
  ram[5320]  = 1;
  ram[5321]  = 1;
  ram[5322]  = 1;
  ram[5323]  = 1;
  ram[5324]  = 1;
  ram[5325]  = 1;
  ram[5326]  = 1;
  ram[5327]  = 1;
  ram[5328]  = 1;
  ram[5329]  = 1;
  ram[5330]  = 1;
  ram[5331]  = 1;
  ram[5332]  = 1;
  ram[5333]  = 1;
  ram[5334]  = 1;
  ram[5335]  = 1;
  ram[5336]  = 1;
  ram[5337]  = 1;
  ram[5338]  = 1;
  ram[5339]  = 1;
  ram[5340]  = 1;
  ram[5341]  = 1;
  ram[5342]  = 1;
  ram[5343]  = 1;
  ram[5344]  = 1;
  ram[5345]  = 1;
  ram[5346]  = 1;
  ram[5347]  = 1;
  ram[5348]  = 1;
  ram[5349]  = 1;
  ram[5350]  = 1;
  ram[5351]  = 1;
  ram[5352]  = 1;
  ram[5353]  = 1;
  ram[5354]  = 1;
  ram[5355]  = 1;
  ram[5356]  = 1;
  ram[5357]  = 1;
  ram[5358]  = 1;
  ram[5359]  = 1;
  ram[5360]  = 1;
  ram[5361]  = 1;
  ram[5362]  = 1;
  ram[5363]  = 1;
  ram[5364]  = 1;
  ram[5365]  = 1;
  ram[5366]  = 1;
  ram[5367]  = 1;
  ram[5368]  = 1;
  ram[5369]  = 1;
  ram[5370]  = 1;
  ram[5371]  = 1;
  ram[5372]  = 1;
  ram[5373]  = 1;
  ram[5374]  = 1;
  ram[5375]  = 1;
  ram[5376]  = 1;
  ram[5377]  = 1;
  ram[5378]  = 1;
  ram[5379]  = 1;
  ram[5380]  = 1;
  ram[5381]  = 1;
  ram[5382]  = 1;
  ram[5383]  = 1;
  ram[5384]  = 1;
  ram[5385]  = 1;
  ram[5386]  = 1;
  ram[5387]  = 1;
  ram[5388]  = 1;
  ram[5389]  = 1;
  ram[5390]  = 1;
  ram[5391]  = 1;
  ram[5392]  = 1;
  ram[5393]  = 1;
  ram[5394]  = 1;
  ram[5395]  = 1;
  ram[5396]  = 1;
  ram[5397]  = 1;
  ram[5398]  = 1;
  ram[5399]  = 1;
  ram[5400]  = 1;
  ram[5401]  = 1;
  ram[5402]  = 1;
  ram[5403]  = 1;
  ram[5404]  = 1;
  ram[5405]  = 1;
  ram[5406]  = 1;
  ram[5407]  = 1;
  ram[5408]  = 1;
  ram[5409]  = 1;
  ram[5410]  = 1;
  ram[5411]  = 1;
  ram[5412]  = 1;
  ram[5413]  = 1;
  ram[5414]  = 1;
  ram[5415]  = 1;
  ram[5416]  = 1;
  ram[5417]  = 1;
  ram[5418]  = 1;
  ram[5419]  = 1;
  ram[5420]  = 1;
  ram[5421]  = 1;
  ram[5422]  = 1;
  ram[5423]  = 1;
  ram[5424]  = 1;
  ram[5425]  = 1;
  ram[5426]  = 1;
  ram[5427]  = 1;
  ram[5428]  = 1;
  ram[5429]  = 1;
  ram[5430]  = 1;
  ram[5431]  = 1;
  ram[5432]  = 1;
  ram[5433]  = 1;
  ram[5434]  = 1;
  ram[5435]  = 1;
  ram[5436]  = 1;
  ram[5437]  = 1;
  ram[5438]  = 1;
  ram[5439]  = 1;
  ram[5440]  = 1;
  ram[5441]  = 1;
  ram[5442]  = 1;
  ram[5443]  = 1;
  ram[5444]  = 1;
  ram[5445]  = 1;
  ram[5446]  = 1;
  ram[5447]  = 1;
  ram[5448]  = 1;
  ram[5449]  = 1;
  ram[5450]  = 1;
  ram[5451]  = 1;
  ram[5452]  = 1;
  ram[5453]  = 1;
  ram[5454]  = 1;
  ram[5455]  = 1;
  ram[5456]  = 1;
  ram[5457]  = 1;
  ram[5458]  = 1;
  ram[5459]  = 1;
  ram[5460]  = 1;
  ram[5461]  = 1;
  ram[5462]  = 1;
  ram[5463]  = 1;
  ram[5464]  = 1;
  ram[5465]  = 1;
  ram[5466]  = 1;
  ram[5467]  = 1;
  ram[5468]  = 1;
  ram[5469]  = 1;
  ram[5470]  = 1;
  ram[5471]  = 1;
  ram[5472]  = 1;
  ram[5473]  = 1;
  ram[5474]  = 1;
  ram[5475]  = 1;
  ram[5476]  = 1;
  ram[5477]  = 1;
  ram[5478]  = 1;
  ram[5479]  = 1;
  ram[5480]  = 1;
  ram[5481]  = 1;
  ram[5482]  = 1;
  ram[5483]  = 1;
  ram[5484]  = 1;
  ram[5485]  = 1;
  ram[5486]  = 1;
  ram[5487]  = 1;
  ram[5488]  = 1;
  ram[5489]  = 1;
  ram[5490]  = 1;
  ram[5491]  = 1;
  ram[5492]  = 1;
  ram[5493]  = 1;
  ram[5494]  = 1;
  ram[5495]  = 1;
  ram[5496]  = 1;
  ram[5497]  = 1;
  ram[5498]  = 1;
  ram[5499]  = 1;
  ram[5500]  = 1;
  ram[5501]  = 1;
  ram[5502]  = 0;
  ram[5503]  = 0;
  ram[5504]  = 0;
  ram[5505]  = 1;
  ram[5506]  = 0;
  ram[5507]  = 0;
  ram[5508]  = 0;
  ram[5509]  = 1;
  ram[5510]  = 1;
  ram[5511]  = 1;
  ram[5512]  = 1;
  ram[5513]  = 1;
  ram[5514]  = 1;
  ram[5515]  = 1;
  ram[5516]  = 1;
  ram[5517]  = 1;
  ram[5518]  = 1;
  ram[5519]  = 1;
  ram[5520]  = 1;
  ram[5521]  = 1;
  ram[5522]  = 1;
  ram[5523]  = 1;
  ram[5524]  = 1;
  ram[5525]  = 1;
  ram[5526]  = 1;
  ram[5527]  = 1;
  ram[5528]  = 1;
  ram[5529]  = 1;
  ram[5530]  = 1;
  ram[5531]  = 1;
  ram[5532]  = 1;
  ram[5533]  = 1;
  ram[5534]  = 1;
  ram[5535]  = 1;
  ram[5536]  = 1;
  ram[5537]  = 1;
  ram[5538]  = 1;
  ram[5539]  = 1;
  ram[5540]  = 1;
  ram[5541]  = 1;
  ram[5542]  = 1;
  ram[5543]  = 1;
  ram[5544]  = 1;
  ram[5545]  = 1;
  ram[5546]  = 1;
  ram[5547]  = 1;
  ram[5548]  = 1;
  ram[5549]  = 1;
  ram[5550]  = 1;
  ram[5551]  = 1;
  ram[5552]  = 1;
  ram[5553]  = 1;
  ram[5554]  = 0;
  ram[5555]  = 0;
  ram[5556]  = 0;
  ram[5557]  = 1;
  ram[5558]  = 1;
  ram[5559]  = 0;
  ram[5560]  = 0;
  ram[5561]  = 0;
  ram[5562]  = 1;
  ram[5563]  = 1;
  ram[5564]  = 1;
  ram[5565]  = 1;
  ram[5566]  = 1;
  ram[5567]  = 1;
  ram[5568]  = 1;
  ram[5569]  = 1;
  ram[5570]  = 1;
  ram[5571]  = 1;
  ram[5572]  = 1;
  ram[5573]  = 1;
  ram[5574]  = 1;
  ram[5575]  = 1;
  ram[5576]  = 1;
  ram[5577]  = 1;
  ram[5578]  = 1;
  ram[5579]  = 1;
  ram[5580]  = 1;
  ram[5581]  = 1;
  ram[5582]  = 1;
  ram[5583]  = 1;
  ram[5584]  = 1;
  ram[5585]  = 1;
  ram[5586]  = 1;
  ram[5587]  = 1;
  ram[5588]  = 1;
  ram[5589]  = 1;
  ram[5590]  = 1;
  ram[5591]  = 0;
  ram[5592]  = 0;
  ram[5593]  = 1;
  ram[5594]  = 1;
  ram[5595]  = 1;
  ram[5596]  = 1;
  ram[5597]  = 1;
  ram[5598]  = 1;
  ram[5599]  = 1;
  ram[5600]  = 1;
  ram[5601]  = 1;
  ram[5602]  = 1;
  ram[5603]  = 1;
  ram[5604]  = 1;
  ram[5605]  = 1;
  ram[5606]  = 1;
  ram[5607]  = 1;
  ram[5608]  = 1;
  ram[5609]  = 1;
  ram[5610]  = 1;
  ram[5611]  = 1;
  ram[5612]  = 1;
  ram[5613]  = 1;
  ram[5614]  = 1;
  ram[5615]  = 1;
  ram[5616]  = 1;
  ram[5617]  = 1;
  ram[5618]  = 1;
  ram[5619]  = 1;
  ram[5620]  = 1;
  ram[5621]  = 1;
  ram[5622]  = 1;
  ram[5623]  = 1;
  ram[5624]  = 1;
  ram[5625]  = 1;
  ram[5626]  = 1;
  ram[5627]  = 1;
  ram[5628]  = 1;
  ram[5629]  = 1;
  ram[5630]  = 1;
  ram[5631]  = 1;
  ram[5632]  = 1;
  ram[5633]  = 1;
  ram[5634]  = 1;
  ram[5635]  = 1;
  ram[5636]  = 1;
  ram[5637]  = 1;
  ram[5638]  = 1;
  ram[5639]  = 1;
  ram[5640]  = 1;
  ram[5641]  = 1;
  ram[5642]  = 1;
  ram[5643]  = 1;
  ram[5644]  = 1;
  ram[5645]  = 1;
  ram[5646]  = 1;
  ram[5647]  = 1;
  ram[5648]  = 1;
  ram[5649]  = 1;
  ram[5650]  = 1;
  ram[5651]  = 1;
  ram[5652]  = 1;
  ram[5653]  = 1;
  ram[5654]  = 1;
  ram[5655]  = 1;
  ram[5656]  = 1;
  ram[5657]  = 1;
  ram[5658]  = 1;
  ram[5659]  = 1;
  ram[5660]  = 1;
  ram[5661]  = 1;
  ram[5662]  = 1;
  ram[5663]  = 1;
  ram[5664]  = 1;
  ram[5665]  = 1;
  ram[5666]  = 1;
  ram[5667]  = 1;
  ram[5668]  = 1;
  ram[5669]  = 1;
  ram[5670]  = 1;
  ram[5671]  = 1;
  ram[5672]  = 1;
  ram[5673]  = 1;
  ram[5674]  = 1;
  ram[5675]  = 1;
  ram[5676]  = 1;
  ram[5677]  = 1;
  ram[5678]  = 1;
  ram[5679]  = 1;
  ram[5680]  = 1;
  ram[5681]  = 1;
  ram[5682]  = 1;
  ram[5683]  = 1;
  ram[5684]  = 1;
  ram[5685]  = 1;
  ram[5686]  = 1;
  ram[5687]  = 1;
  ram[5688]  = 1;
  ram[5689]  = 1;
  ram[5690]  = 1;
  ram[5691]  = 1;
  ram[5692]  = 1;
  ram[5693]  = 1;
  ram[5694]  = 1;
  ram[5695]  = 1;
  ram[5696]  = 1;
  ram[5697]  = 1;
  ram[5698]  = 1;
  ram[5699]  = 1;
  ram[5700]  = 1;
  ram[5701]  = 1;
  ram[5702]  = 1;
  ram[5703]  = 1;
  ram[5704]  = 1;
  ram[5705]  = 1;
  ram[5706]  = 1;
  ram[5707]  = 1;
  ram[5708]  = 1;
  ram[5709]  = 1;
  ram[5710]  = 1;
  ram[5711]  = 1;
  ram[5712]  = 1;
  ram[5713]  = 1;
  ram[5714]  = 1;
  ram[5715]  = 1;
  ram[5716]  = 1;
  ram[5717]  = 1;
  ram[5718]  = 1;
  ram[5719]  = 1;
  ram[5720]  = 1;
  ram[5721]  = 1;
  ram[5722]  = 1;
  ram[5723]  = 1;
  ram[5724]  = 1;
  ram[5725]  = 1;
  ram[5726]  = 1;
  ram[5727]  = 1;
  ram[5728]  = 1;
  ram[5729]  = 1;
  ram[5730]  = 1;
  ram[5731]  = 1;
  ram[5732]  = 1;
  ram[5733]  = 1;
  ram[5734]  = 1;
  ram[5735]  = 1;
  ram[5736]  = 1;
  ram[5737]  = 1;
  ram[5738]  = 1;
  ram[5739]  = 1;
  ram[5740]  = 1;
  ram[5741]  = 1;
  ram[5742]  = 1;
  ram[5743]  = 1;
  ram[5744]  = 1;
  ram[5745]  = 1;
  ram[5746]  = 1;
  ram[5747]  = 1;
  ram[5748]  = 1;
  ram[5749]  = 1;
  ram[5750]  = 1;
  ram[5751]  = 1;
  ram[5752]  = 1;
  ram[5753]  = 1;
  ram[5754]  = 1;
  ram[5755]  = 1;
  ram[5756]  = 1;
  ram[5757]  = 1;
  ram[5758]  = 1;
  ram[5759]  = 1;
  ram[5760]  = 1;
  ram[5761]  = 1;
  ram[5762]  = 1;
  ram[5763]  = 1;
  ram[5764]  = 1;
  ram[5765]  = 1;
  ram[5766]  = 1;
  ram[5767]  = 1;
  ram[5768]  = 1;
  ram[5769]  = 1;
  ram[5770]  = 1;
  ram[5771]  = 1;
  ram[5772]  = 1;
  ram[5773]  = 1;
  ram[5774]  = 1;
  ram[5775]  = 1;
  ram[5776]  = 1;
  ram[5777]  = 1;
  ram[5778]  = 1;
  ram[5779]  = 1;
  ram[5780]  = 1;
  ram[5781]  = 1;
  ram[5782]  = 1;
  ram[5783]  = 1;
  ram[5784]  = 1;
  ram[5785]  = 1;
  ram[5786]  = 1;
  ram[5787]  = 1;
  ram[5788]  = 1;
  ram[5789]  = 1;
  ram[5790]  = 1;
  ram[5791]  = 1;
  ram[5792]  = 1;
  ram[5793]  = 1;
  ram[5794]  = 1;
  ram[5795]  = 1;
  ram[5796]  = 1;
  ram[5797]  = 1;
  ram[5798]  = 1;
  ram[5799]  = 1;
  ram[5800]  = 1;
  ram[5801]  = 0;
  ram[5802]  = 0;
  ram[5803]  = 1;
  ram[5804]  = 1;
  ram[5805]  = 1;
  ram[5806]  = 1;
  ram[5807]  = 1;
  ram[5808]  = 0;
  ram[5809]  = 0;
  ram[5810]  = 1;
  ram[5811]  = 1;
  ram[5812]  = 1;
  ram[5813]  = 1;
  ram[5814]  = 1;
  ram[5815]  = 1;
  ram[5816]  = 1;
  ram[5817]  = 1;
  ram[5818]  = 1;
  ram[5819]  = 1;
  ram[5820]  = 1;
  ram[5821]  = 1;
  ram[5822]  = 1;
  ram[5823]  = 1;
  ram[5824]  = 1;
  ram[5825]  = 1;
  ram[5826]  = 1;
  ram[5827]  = 1;
  ram[5828]  = 1;
  ram[5829]  = 1;
  ram[5830]  = 1;
  ram[5831]  = 1;
  ram[5832]  = 1;
  ram[5833]  = 1;
  ram[5834]  = 1;
  ram[5835]  = 1;
  ram[5836]  = 1;
  ram[5837]  = 1;
  ram[5838]  = 1;
  ram[5839]  = 1;
  ram[5840]  = 1;
  ram[5841]  = 1;
  ram[5842]  = 1;
  ram[5843]  = 1;
  ram[5844]  = 1;
  ram[5845]  = 1;
  ram[5846]  = 1;
  ram[5847]  = 1;
  ram[5848]  = 1;
  ram[5849]  = 1;
  ram[5850]  = 1;
  ram[5851]  = 1;
  ram[5852]  = 1;
  ram[5853]  = 1;
  ram[5854]  = 0;
  ram[5855]  = 0;
  ram[5856]  = 1;
  ram[5857]  = 1;
  ram[5858]  = 1;
  ram[5859]  = 1;
  ram[5860]  = 1;
  ram[5861]  = 0;
  ram[5862]  = 1;
  ram[5863]  = 1;
  ram[5864]  = 1;
  ram[5865]  = 1;
  ram[5866]  = 1;
  ram[5867]  = 1;
  ram[5868]  = 1;
  ram[5869]  = 1;
  ram[5870]  = 1;
  ram[5871]  = 1;
  ram[5872]  = 1;
  ram[5873]  = 1;
  ram[5874]  = 1;
  ram[5875]  = 1;
  ram[5876]  = 1;
  ram[5877]  = 1;
  ram[5878]  = 1;
  ram[5879]  = 1;
  ram[5880]  = 1;
  ram[5881]  = 1;
  ram[5882]  = 1;
  ram[5883]  = 1;
  ram[5884]  = 1;
  ram[5885]  = 1;
  ram[5886]  = 1;
  ram[5887]  = 1;
  ram[5888]  = 1;
  ram[5889]  = 1;
  ram[5890]  = 1;
  ram[5891]  = 0;
  ram[5892]  = 0;
  ram[5893]  = 1;
  ram[5894]  = 1;
  ram[5895]  = 1;
  ram[5896]  = 1;
  ram[5897]  = 1;
  ram[5898]  = 1;
  ram[5899]  = 1;
  ram[5900]  = 1;
  ram[5901]  = 1;
  ram[5902]  = 1;
  ram[5903]  = 1;
  ram[5904]  = 1;
  ram[5905]  = 1;
  ram[5906]  = 1;
  ram[5907]  = 1;
  ram[5908]  = 1;
  ram[5909]  = 1;
  ram[5910]  = 1;
  ram[5911]  = 1;
  ram[5912]  = 1;
  ram[5913]  = 1;
  ram[5914]  = 1;
  ram[5915]  = 1;
  ram[5916]  = 1;
  ram[5917]  = 1;
  ram[5918]  = 1;
  ram[5919]  = 1;
  ram[5920]  = 1;
  ram[5921]  = 1;
  ram[5922]  = 1;
  ram[5923]  = 1;
  ram[5924]  = 1;
  ram[5925]  = 1;
  ram[5926]  = 1;
  ram[5927]  = 1;
  ram[5928]  = 1;
  ram[5929]  = 1;
  ram[5930]  = 1;
  ram[5931]  = 1;
  ram[5932]  = 1;
  ram[5933]  = 1;
  ram[5934]  = 1;
  ram[5935]  = 1;
  ram[5936]  = 1;
  ram[5937]  = 1;
  ram[5938]  = 1;
  ram[5939]  = 1;
  ram[5940]  = 1;
  ram[5941]  = 1;
  ram[5942]  = 1;
  ram[5943]  = 1;
  ram[5944]  = 1;
  ram[5945]  = 1;
  ram[5946]  = 1;
  ram[5947]  = 1;
  ram[5948]  = 1;
  ram[5949]  = 1;
  ram[5950]  = 1;
  ram[5951]  = 1;
  ram[5952]  = 1;
  ram[5953]  = 1;
  ram[5954]  = 1;
  ram[5955]  = 1;
  ram[5956]  = 1;
  ram[5957]  = 1;
  ram[5958]  = 1;
  ram[5959]  = 1;
  ram[5960]  = 1;
  ram[5961]  = 1;
  ram[5962]  = 1;
  ram[5963]  = 1;
  ram[5964]  = 1;
  ram[5965]  = 1;
  ram[5966]  = 1;
  ram[5967]  = 1;
  ram[5968]  = 1;
  ram[5969]  = 1;
  ram[5970]  = 1;
  ram[5971]  = 1;
  ram[5972]  = 1;
  ram[5973]  = 1;
  ram[5974]  = 1;
  ram[5975]  = 1;
  ram[5976]  = 1;
  ram[5977]  = 1;
  ram[5978]  = 1;
  ram[5979]  = 1;
  ram[5980]  = 1;
  ram[5981]  = 1;
  ram[5982]  = 1;
  ram[5983]  = 1;
  ram[5984]  = 1;
  ram[5985]  = 1;
  ram[5986]  = 1;
  ram[5987]  = 1;
  ram[5988]  = 1;
  ram[5989]  = 1;
  ram[5990]  = 1;
  ram[5991]  = 1;
  ram[5992]  = 1;
  ram[5993]  = 1;
  ram[5994]  = 1;
  ram[5995]  = 1;
  ram[5996]  = 1;
  ram[5997]  = 1;
  ram[5998]  = 1;
  ram[5999]  = 1;
  ram[6000]  = 1;
  ram[6001]  = 1;
  ram[6002]  = 1;
  ram[6003]  = 1;
  ram[6004]  = 1;
  ram[6005]  = 1;
  ram[6006]  = 1;
  ram[6007]  = 1;
  ram[6008]  = 1;
  ram[6009]  = 1;
  ram[6010]  = 1;
  ram[6011]  = 1;
  ram[6012]  = 1;
  ram[6013]  = 1;
  ram[6014]  = 1;
  ram[6015]  = 1;
  ram[6016]  = 1;
  ram[6017]  = 1;
  ram[6018]  = 1;
  ram[6019]  = 1;
  ram[6020]  = 1;
  ram[6021]  = 1;
  ram[6022]  = 1;
  ram[6023]  = 1;
  ram[6024]  = 1;
  ram[6025]  = 1;
  ram[6026]  = 1;
  ram[6027]  = 1;
  ram[6028]  = 1;
  ram[6029]  = 1;
  ram[6030]  = 1;
  ram[6031]  = 1;
  ram[6032]  = 1;
  ram[6033]  = 1;
  ram[6034]  = 1;
  ram[6035]  = 1;
  ram[6036]  = 1;
  ram[6037]  = 1;
  ram[6038]  = 1;
  ram[6039]  = 1;
  ram[6040]  = 1;
  ram[6041]  = 1;
  ram[6042]  = 1;
  ram[6043]  = 1;
  ram[6044]  = 1;
  ram[6045]  = 1;
  ram[6046]  = 1;
  ram[6047]  = 1;
  ram[6048]  = 1;
  ram[6049]  = 1;
  ram[6050]  = 1;
  ram[6051]  = 1;
  ram[6052]  = 1;
  ram[6053]  = 1;
  ram[6054]  = 1;
  ram[6055]  = 1;
  ram[6056]  = 1;
  ram[6057]  = 1;
  ram[6058]  = 1;
  ram[6059]  = 1;
  ram[6060]  = 1;
  ram[6061]  = 1;
  ram[6062]  = 1;
  ram[6063]  = 1;
  ram[6064]  = 1;
  ram[6065]  = 1;
  ram[6066]  = 1;
  ram[6067]  = 1;
  ram[6068]  = 1;
  ram[6069]  = 1;
  ram[6070]  = 1;
  ram[6071]  = 1;
  ram[6072]  = 1;
  ram[6073]  = 1;
  ram[6074]  = 1;
  ram[6075]  = 1;
  ram[6076]  = 1;
  ram[6077]  = 1;
  ram[6078]  = 1;
  ram[6079]  = 1;
  ram[6080]  = 1;
  ram[6081]  = 1;
  ram[6082]  = 1;
  ram[6083]  = 1;
  ram[6084]  = 1;
  ram[6085]  = 1;
  ram[6086]  = 1;
  ram[6087]  = 1;
  ram[6088]  = 1;
  ram[6089]  = 1;
  ram[6090]  = 1;
  ram[6091]  = 1;
  ram[6092]  = 1;
  ram[6093]  = 1;
  ram[6094]  = 1;
  ram[6095]  = 1;
  ram[6096]  = 1;
  ram[6097]  = 1;
  ram[6098]  = 1;
  ram[6099]  = 1;
  ram[6100]  = 1;
  ram[6101]  = 0;
  ram[6102]  = 0;
  ram[6103]  = 1;
  ram[6104]  = 1;
  ram[6105]  = 1;
  ram[6106]  = 1;
  ram[6107]  = 1;
  ram[6108]  = 0;
  ram[6109]  = 0;
  ram[6110]  = 1;
  ram[6111]  = 1;
  ram[6112]  = 1;
  ram[6113]  = 1;
  ram[6114]  = 1;
  ram[6115]  = 1;
  ram[6116]  = 1;
  ram[6117]  = 1;
  ram[6118]  = 1;
  ram[6119]  = 1;
  ram[6120]  = 1;
  ram[6121]  = 1;
  ram[6122]  = 1;
  ram[6123]  = 1;
  ram[6124]  = 1;
  ram[6125]  = 1;
  ram[6126]  = 1;
  ram[6127]  = 1;
  ram[6128]  = 1;
  ram[6129]  = 1;
  ram[6130]  = 1;
  ram[6131]  = 1;
  ram[6132]  = 1;
  ram[6133]  = 1;
  ram[6134]  = 1;
  ram[6135]  = 1;
  ram[6136]  = 1;
  ram[6137]  = 1;
  ram[6138]  = 1;
  ram[6139]  = 1;
  ram[6140]  = 1;
  ram[6141]  = 1;
  ram[6142]  = 1;
  ram[6143]  = 1;
  ram[6144]  = 1;
  ram[6145]  = 1;
  ram[6146]  = 1;
  ram[6147]  = 1;
  ram[6148]  = 1;
  ram[6149]  = 1;
  ram[6150]  = 1;
  ram[6151]  = 1;
  ram[6152]  = 1;
  ram[6153]  = 0;
  ram[6154]  = 0;
  ram[6155]  = 1;
  ram[6156]  = 1;
  ram[6157]  = 1;
  ram[6158]  = 1;
  ram[6159]  = 1;
  ram[6160]  = 1;
  ram[6161]  = 0;
  ram[6162]  = 0;
  ram[6163]  = 1;
  ram[6164]  = 1;
  ram[6165]  = 1;
  ram[6166]  = 1;
  ram[6167]  = 1;
  ram[6168]  = 1;
  ram[6169]  = 1;
  ram[6170]  = 1;
  ram[6171]  = 1;
  ram[6172]  = 1;
  ram[6173]  = 1;
  ram[6174]  = 1;
  ram[6175]  = 1;
  ram[6176]  = 1;
  ram[6177]  = 1;
  ram[6178]  = 1;
  ram[6179]  = 1;
  ram[6180]  = 1;
  ram[6181]  = 1;
  ram[6182]  = 1;
  ram[6183]  = 1;
  ram[6184]  = 1;
  ram[6185]  = 1;
  ram[6186]  = 1;
  ram[6187]  = 1;
  ram[6188]  = 1;
  ram[6189]  = 1;
  ram[6190]  = 1;
  ram[6191]  = 0;
  ram[6192]  = 0;
  ram[6193]  = 1;
  ram[6194]  = 1;
  ram[6195]  = 1;
  ram[6196]  = 1;
  ram[6197]  = 1;
  ram[6198]  = 1;
  ram[6199]  = 1;
  ram[6200]  = 1;
  ram[6201]  = 1;
  ram[6202]  = 1;
  ram[6203]  = 1;
  ram[6204]  = 1;
  ram[6205]  = 1;
  ram[6206]  = 1;
  ram[6207]  = 1;
  ram[6208]  = 1;
  ram[6209]  = 1;
  ram[6210]  = 1;
  ram[6211]  = 1;
  ram[6212]  = 1;
  ram[6213]  = 1;
  ram[6214]  = 1;
  ram[6215]  = 1;
  ram[6216]  = 1;
  ram[6217]  = 1;
  ram[6218]  = 1;
  ram[6219]  = 1;
  ram[6220]  = 1;
  ram[6221]  = 1;
  ram[6222]  = 1;
  ram[6223]  = 1;
  ram[6224]  = 1;
  ram[6225]  = 1;
  ram[6226]  = 1;
  ram[6227]  = 1;
  ram[6228]  = 1;
  ram[6229]  = 1;
  ram[6230]  = 1;
  ram[6231]  = 1;
  ram[6232]  = 1;
  ram[6233]  = 1;
  ram[6234]  = 1;
  ram[6235]  = 1;
  ram[6236]  = 1;
  ram[6237]  = 1;
  ram[6238]  = 1;
  ram[6239]  = 1;
  ram[6240]  = 1;
  ram[6241]  = 1;
  ram[6242]  = 1;
  ram[6243]  = 1;
  ram[6244]  = 1;
  ram[6245]  = 1;
  ram[6246]  = 1;
  ram[6247]  = 1;
  ram[6248]  = 1;
  ram[6249]  = 1;
  ram[6250]  = 1;
  ram[6251]  = 1;
  ram[6252]  = 1;
  ram[6253]  = 1;
  ram[6254]  = 1;
  ram[6255]  = 1;
  ram[6256]  = 1;
  ram[6257]  = 1;
  ram[6258]  = 1;
  ram[6259]  = 1;
  ram[6260]  = 1;
  ram[6261]  = 1;
  ram[6262]  = 1;
  ram[6263]  = 1;
  ram[6264]  = 1;
  ram[6265]  = 1;
  ram[6266]  = 1;
  ram[6267]  = 1;
  ram[6268]  = 1;
  ram[6269]  = 1;
  ram[6270]  = 1;
  ram[6271]  = 1;
  ram[6272]  = 1;
  ram[6273]  = 1;
  ram[6274]  = 1;
  ram[6275]  = 1;
  ram[6276]  = 1;
  ram[6277]  = 1;
  ram[6278]  = 1;
  ram[6279]  = 1;
  ram[6280]  = 1;
  ram[6281]  = 1;
  ram[6282]  = 1;
  ram[6283]  = 1;
  ram[6284]  = 1;
  ram[6285]  = 1;
  ram[6286]  = 1;
  ram[6287]  = 1;
  ram[6288]  = 1;
  ram[6289]  = 1;
  ram[6290]  = 1;
  ram[6291]  = 1;
  ram[6292]  = 1;
  ram[6293]  = 1;
  ram[6294]  = 1;
  ram[6295]  = 1;
  ram[6296]  = 1;
  ram[6297]  = 1;
  ram[6298]  = 1;
  ram[6299]  = 1;
  ram[6300]  = 1;
  ram[6301]  = 1;
  ram[6302]  = 1;
  ram[6303]  = 1;
  ram[6304]  = 1;
  ram[6305]  = 1;
  ram[6306]  = 1;
  ram[6307]  = 1;
  ram[6308]  = 1;
  ram[6309]  = 1;
  ram[6310]  = 1;
  ram[6311]  = 1;
  ram[6312]  = 1;
  ram[6313]  = 1;
  ram[6314]  = 1;
  ram[6315]  = 1;
  ram[6316]  = 1;
  ram[6317]  = 1;
  ram[6318]  = 1;
  ram[6319]  = 1;
  ram[6320]  = 1;
  ram[6321]  = 1;
  ram[6322]  = 1;
  ram[6323]  = 1;
  ram[6324]  = 1;
  ram[6325]  = 1;
  ram[6326]  = 1;
  ram[6327]  = 1;
  ram[6328]  = 1;
  ram[6329]  = 1;
  ram[6330]  = 1;
  ram[6331]  = 1;
  ram[6332]  = 1;
  ram[6333]  = 1;
  ram[6334]  = 1;
  ram[6335]  = 1;
  ram[6336]  = 1;
  ram[6337]  = 1;
  ram[6338]  = 1;
  ram[6339]  = 1;
  ram[6340]  = 1;
  ram[6341]  = 1;
  ram[6342]  = 1;
  ram[6343]  = 1;
  ram[6344]  = 1;
  ram[6345]  = 1;
  ram[6346]  = 1;
  ram[6347]  = 1;
  ram[6348]  = 1;
  ram[6349]  = 1;
  ram[6350]  = 1;
  ram[6351]  = 1;
  ram[6352]  = 1;
  ram[6353]  = 1;
  ram[6354]  = 1;
  ram[6355]  = 1;
  ram[6356]  = 1;
  ram[6357]  = 1;
  ram[6358]  = 1;
  ram[6359]  = 1;
  ram[6360]  = 1;
  ram[6361]  = 1;
  ram[6362]  = 1;
  ram[6363]  = 1;
  ram[6364]  = 1;
  ram[6365]  = 1;
  ram[6366]  = 1;
  ram[6367]  = 1;
  ram[6368]  = 1;
  ram[6369]  = 1;
  ram[6370]  = 1;
  ram[6371]  = 1;
  ram[6372]  = 1;
  ram[6373]  = 1;
  ram[6374]  = 1;
  ram[6375]  = 1;
  ram[6376]  = 1;
  ram[6377]  = 1;
  ram[6378]  = 1;
  ram[6379]  = 1;
  ram[6380]  = 1;
  ram[6381]  = 1;
  ram[6382]  = 1;
  ram[6383]  = 1;
  ram[6384]  = 1;
  ram[6385]  = 1;
  ram[6386]  = 1;
  ram[6387]  = 1;
  ram[6388]  = 1;
  ram[6389]  = 1;
  ram[6390]  = 1;
  ram[6391]  = 1;
  ram[6392]  = 1;
  ram[6393]  = 1;
  ram[6394]  = 1;
  ram[6395]  = 1;
  ram[6396]  = 1;
  ram[6397]  = 1;
  ram[6398]  = 1;
  ram[6399]  = 1;
  ram[6400]  = 1;
  ram[6401]  = 0;
  ram[6402]  = 1;
  ram[6403]  = 1;
  ram[6404]  = 1;
  ram[6405]  = 1;
  ram[6406]  = 1;
  ram[6407]  = 1;
  ram[6408]  = 1;
  ram[6409]  = 0;
  ram[6410]  = 1;
  ram[6411]  = 1;
  ram[6412]  = 1;
  ram[6413]  = 1;
  ram[6414]  = 1;
  ram[6415]  = 1;
  ram[6416]  = 1;
  ram[6417]  = 1;
  ram[6418]  = 1;
  ram[6419]  = 1;
  ram[6420]  = 1;
  ram[6421]  = 1;
  ram[6422]  = 1;
  ram[6423]  = 1;
  ram[6424]  = 1;
  ram[6425]  = 1;
  ram[6426]  = 1;
  ram[6427]  = 1;
  ram[6428]  = 1;
  ram[6429]  = 1;
  ram[6430]  = 1;
  ram[6431]  = 1;
  ram[6432]  = 1;
  ram[6433]  = 1;
  ram[6434]  = 1;
  ram[6435]  = 1;
  ram[6436]  = 1;
  ram[6437]  = 1;
  ram[6438]  = 1;
  ram[6439]  = 1;
  ram[6440]  = 1;
  ram[6441]  = 1;
  ram[6442]  = 1;
  ram[6443]  = 1;
  ram[6444]  = 1;
  ram[6445]  = 1;
  ram[6446]  = 1;
  ram[6447]  = 1;
  ram[6448]  = 1;
  ram[6449]  = 1;
  ram[6450]  = 1;
  ram[6451]  = 1;
  ram[6452]  = 1;
  ram[6453]  = 0;
  ram[6454]  = 1;
  ram[6455]  = 1;
  ram[6456]  = 1;
  ram[6457]  = 1;
  ram[6458]  = 1;
  ram[6459]  = 1;
  ram[6460]  = 1;
  ram[6461]  = 1;
  ram[6462]  = 0;
  ram[6463]  = 1;
  ram[6464]  = 1;
  ram[6465]  = 1;
  ram[6466]  = 1;
  ram[6467]  = 1;
  ram[6468]  = 1;
  ram[6469]  = 1;
  ram[6470]  = 1;
  ram[6471]  = 1;
  ram[6472]  = 1;
  ram[6473]  = 1;
  ram[6474]  = 1;
  ram[6475]  = 1;
  ram[6476]  = 1;
  ram[6477]  = 1;
  ram[6478]  = 1;
  ram[6479]  = 1;
  ram[6480]  = 1;
  ram[6481]  = 1;
  ram[6482]  = 1;
  ram[6483]  = 1;
  ram[6484]  = 1;
  ram[6485]  = 1;
  ram[6486]  = 1;
  ram[6487]  = 1;
  ram[6488]  = 1;
  ram[6489]  = 1;
  ram[6490]  = 1;
  ram[6491]  = 0;
  ram[6492]  = 0;
  ram[6493]  = 1;
  ram[6494]  = 1;
  ram[6495]  = 1;
  ram[6496]  = 1;
  ram[6497]  = 1;
  ram[6498]  = 1;
  ram[6499]  = 1;
  ram[6500]  = 1;
  ram[6501]  = 1;
  ram[6502]  = 1;
  ram[6503]  = 1;
  ram[6504]  = 1;
  ram[6505]  = 1;
  ram[6506]  = 1;
  ram[6507]  = 1;
  ram[6508]  = 1;
  ram[6509]  = 1;
  ram[6510]  = 1;
  ram[6511]  = 1;
  ram[6512]  = 1;
  ram[6513]  = 1;
  ram[6514]  = 1;
  ram[6515]  = 1;
  ram[6516]  = 1;
  ram[6517]  = 1;
  ram[6518]  = 1;
  ram[6519]  = 1;
  ram[6520]  = 1;
  ram[6521]  = 1;
  ram[6522]  = 1;
  ram[6523]  = 1;
  ram[6524]  = 1;
  ram[6525]  = 1;
  ram[6526]  = 1;
  ram[6527]  = 1;
  ram[6528]  = 1;
  ram[6529]  = 1;
  ram[6530]  = 1;
  ram[6531]  = 1;
  ram[6532]  = 1;
  ram[6533]  = 1;
  ram[6534]  = 1;
  ram[6535]  = 1;
  ram[6536]  = 1;
  ram[6537]  = 1;
  ram[6538]  = 1;
  ram[6539]  = 1;
  ram[6540]  = 1;
  ram[6541]  = 1;
  ram[6542]  = 1;
  ram[6543]  = 1;
  ram[6544]  = 1;
  ram[6545]  = 1;
  ram[6546]  = 1;
  ram[6547]  = 1;
  ram[6548]  = 1;
  ram[6549]  = 1;
  ram[6550]  = 1;
  ram[6551]  = 1;
  ram[6552]  = 1;
  ram[6553]  = 1;
  ram[6554]  = 1;
  ram[6555]  = 1;
  ram[6556]  = 1;
  ram[6557]  = 1;
  ram[6558]  = 1;
  ram[6559]  = 1;
  ram[6560]  = 1;
  ram[6561]  = 1;
  ram[6562]  = 1;
  ram[6563]  = 1;
  ram[6564]  = 1;
  ram[6565]  = 1;
  ram[6566]  = 1;
  ram[6567]  = 1;
  ram[6568]  = 1;
  ram[6569]  = 1;
  ram[6570]  = 1;
  ram[6571]  = 1;
  ram[6572]  = 1;
  ram[6573]  = 1;
  ram[6574]  = 1;
  ram[6575]  = 1;
  ram[6576]  = 1;
  ram[6577]  = 1;
  ram[6578]  = 1;
  ram[6579]  = 1;
  ram[6580]  = 1;
  ram[6581]  = 1;
  ram[6582]  = 1;
  ram[6583]  = 1;
  ram[6584]  = 1;
  ram[6585]  = 1;
  ram[6586]  = 1;
  ram[6587]  = 1;
  ram[6588]  = 1;
  ram[6589]  = 1;
  ram[6590]  = 1;
  ram[6591]  = 1;
  ram[6592]  = 1;
  ram[6593]  = 1;
  ram[6594]  = 1;
  ram[6595]  = 1;
  ram[6596]  = 1;
  ram[6597]  = 1;
  ram[6598]  = 1;
  ram[6599]  = 1;
  ram[6600]  = 1;
  ram[6601]  = 1;
  ram[6602]  = 1;
  ram[6603]  = 1;
  ram[6604]  = 1;
  ram[6605]  = 1;
  ram[6606]  = 1;
  ram[6607]  = 1;
  ram[6608]  = 1;
  ram[6609]  = 1;
  ram[6610]  = 1;
  ram[6611]  = 1;
  ram[6612]  = 1;
  ram[6613]  = 1;
  ram[6614]  = 1;
  ram[6615]  = 1;
  ram[6616]  = 1;
  ram[6617]  = 1;
  ram[6618]  = 1;
  ram[6619]  = 1;
  ram[6620]  = 1;
  ram[6621]  = 1;
  ram[6622]  = 1;
  ram[6623]  = 1;
  ram[6624]  = 1;
  ram[6625]  = 1;
  ram[6626]  = 1;
  ram[6627]  = 1;
  ram[6628]  = 1;
  ram[6629]  = 1;
  ram[6630]  = 1;
  ram[6631]  = 1;
  ram[6632]  = 1;
  ram[6633]  = 1;
  ram[6634]  = 1;
  ram[6635]  = 1;
  ram[6636]  = 1;
  ram[6637]  = 1;
  ram[6638]  = 1;
  ram[6639]  = 1;
  ram[6640]  = 1;
  ram[6641]  = 1;
  ram[6642]  = 1;
  ram[6643]  = 1;
  ram[6644]  = 1;
  ram[6645]  = 1;
  ram[6646]  = 1;
  ram[6647]  = 1;
  ram[6648]  = 1;
  ram[6649]  = 1;
  ram[6650]  = 1;
  ram[6651]  = 1;
  ram[6652]  = 1;
  ram[6653]  = 1;
  ram[6654]  = 1;
  ram[6655]  = 1;
  ram[6656]  = 1;
  ram[6657]  = 1;
  ram[6658]  = 1;
  ram[6659]  = 1;
  ram[6660]  = 1;
  ram[6661]  = 1;
  ram[6662]  = 1;
  ram[6663]  = 1;
  ram[6664]  = 1;
  ram[6665]  = 1;
  ram[6666]  = 1;
  ram[6667]  = 1;
  ram[6668]  = 1;
  ram[6669]  = 1;
  ram[6670]  = 1;
  ram[6671]  = 1;
  ram[6672]  = 1;
  ram[6673]  = 1;
  ram[6674]  = 1;
  ram[6675]  = 1;
  ram[6676]  = 1;
  ram[6677]  = 1;
  ram[6678]  = 1;
  ram[6679]  = 1;
  ram[6680]  = 1;
  ram[6681]  = 1;
  ram[6682]  = 1;
  ram[6683]  = 1;
  ram[6684]  = 1;
  ram[6685]  = 1;
  ram[6686]  = 1;
  ram[6687]  = 1;
  ram[6688]  = 1;
  ram[6689]  = 1;
  ram[6690]  = 1;
  ram[6691]  = 1;
  ram[6692]  = 1;
  ram[6693]  = 1;
  ram[6694]  = 1;
  ram[6695]  = 1;
  ram[6696]  = 1;
  ram[6697]  = 1;
  ram[6698]  = 1;
  ram[6699]  = 1;
  ram[6700]  = 0;
  ram[6701]  = 0;
  ram[6702]  = 1;
  ram[6703]  = 1;
  ram[6704]  = 1;
  ram[6705]  = 1;
  ram[6706]  = 1;
  ram[6707]  = 1;
  ram[6708]  = 1;
  ram[6709]  = 1;
  ram[6710]  = 1;
  ram[6711]  = 1;
  ram[6712]  = 1;
  ram[6713]  = 1;
  ram[6714]  = 1;
  ram[6715]  = 1;
  ram[6716]  = 1;
  ram[6717]  = 1;
  ram[6718]  = 1;
  ram[6719]  = 1;
  ram[6720]  = 1;
  ram[6721]  = 1;
  ram[6722]  = 1;
  ram[6723]  = 1;
  ram[6724]  = 1;
  ram[6725]  = 1;
  ram[6726]  = 1;
  ram[6727]  = 1;
  ram[6728]  = 1;
  ram[6729]  = 1;
  ram[6730]  = 1;
  ram[6731]  = 1;
  ram[6732]  = 1;
  ram[6733]  = 1;
  ram[6734]  = 1;
  ram[6735]  = 1;
  ram[6736]  = 1;
  ram[6737]  = 1;
  ram[6738]  = 1;
  ram[6739]  = 1;
  ram[6740]  = 1;
  ram[6741]  = 1;
  ram[6742]  = 1;
  ram[6743]  = 1;
  ram[6744]  = 1;
  ram[6745]  = 1;
  ram[6746]  = 1;
  ram[6747]  = 1;
  ram[6748]  = 1;
  ram[6749]  = 1;
  ram[6750]  = 1;
  ram[6751]  = 1;
  ram[6752]  = 1;
  ram[6753]  = 0;
  ram[6754]  = 1;
  ram[6755]  = 1;
  ram[6756]  = 1;
  ram[6757]  = 1;
  ram[6758]  = 1;
  ram[6759]  = 1;
  ram[6760]  = 1;
  ram[6761]  = 1;
  ram[6762]  = 0;
  ram[6763]  = 0;
  ram[6764]  = 1;
  ram[6765]  = 1;
  ram[6766]  = 1;
  ram[6767]  = 1;
  ram[6768]  = 1;
  ram[6769]  = 1;
  ram[6770]  = 1;
  ram[6771]  = 1;
  ram[6772]  = 1;
  ram[6773]  = 1;
  ram[6774]  = 1;
  ram[6775]  = 1;
  ram[6776]  = 1;
  ram[6777]  = 1;
  ram[6778]  = 1;
  ram[6779]  = 1;
  ram[6780]  = 1;
  ram[6781]  = 1;
  ram[6782]  = 1;
  ram[6783]  = 1;
  ram[6784]  = 1;
  ram[6785]  = 1;
  ram[6786]  = 1;
  ram[6787]  = 1;
  ram[6788]  = 1;
  ram[6789]  = 1;
  ram[6790]  = 1;
  ram[6791]  = 0;
  ram[6792]  = 0;
  ram[6793]  = 1;
  ram[6794]  = 1;
  ram[6795]  = 1;
  ram[6796]  = 1;
  ram[6797]  = 1;
  ram[6798]  = 1;
  ram[6799]  = 1;
  ram[6800]  = 1;
  ram[6801]  = 1;
  ram[6802]  = 1;
  ram[6803]  = 1;
  ram[6804]  = 1;
  ram[6805]  = 1;
  ram[6806]  = 1;
  ram[6807]  = 1;
  ram[6808]  = 1;
  ram[6809]  = 1;
  ram[6810]  = 1;
  ram[6811]  = 1;
  ram[6812]  = 1;
  ram[6813]  = 1;
  ram[6814]  = 1;
  ram[6815]  = 1;
  ram[6816]  = 1;
  ram[6817]  = 1;
  ram[6818]  = 1;
  ram[6819]  = 1;
  ram[6820]  = 1;
  ram[6821]  = 1;
  ram[6822]  = 1;
  ram[6823]  = 1;
  ram[6824]  = 1;
  ram[6825]  = 1;
  ram[6826]  = 1;
  ram[6827]  = 1;
  ram[6828]  = 1;
  ram[6829]  = 1;
  ram[6830]  = 1;
  ram[6831]  = 1;
  ram[6832]  = 1;
  ram[6833]  = 1;
  ram[6834]  = 1;
  ram[6835]  = 1;
  ram[6836]  = 1;
  ram[6837]  = 1;
  ram[6838]  = 1;
  ram[6839]  = 1;
  ram[6840]  = 1;
  ram[6841]  = 1;
  ram[6842]  = 1;
  ram[6843]  = 1;
  ram[6844]  = 1;
  ram[6845]  = 1;
  ram[6846]  = 1;
  ram[6847]  = 1;
  ram[6848]  = 1;
  ram[6849]  = 1;
  ram[6850]  = 1;
  ram[6851]  = 1;
  ram[6852]  = 1;
  ram[6853]  = 1;
  ram[6854]  = 1;
  ram[6855]  = 1;
  ram[6856]  = 1;
  ram[6857]  = 1;
  ram[6858]  = 1;
  ram[6859]  = 1;
  ram[6860]  = 1;
  ram[6861]  = 1;
  ram[6862]  = 1;
  ram[6863]  = 1;
  ram[6864]  = 1;
  ram[6865]  = 1;
  ram[6866]  = 1;
  ram[6867]  = 1;
  ram[6868]  = 1;
  ram[6869]  = 1;
  ram[6870]  = 1;
  ram[6871]  = 1;
  ram[6872]  = 1;
  ram[6873]  = 1;
  ram[6874]  = 1;
  ram[6875]  = 1;
  ram[6876]  = 1;
  ram[6877]  = 1;
  ram[6878]  = 1;
  ram[6879]  = 1;
  ram[6880]  = 1;
  ram[6881]  = 1;
  ram[6882]  = 1;
  ram[6883]  = 1;
  ram[6884]  = 1;
  ram[6885]  = 1;
  ram[6886]  = 1;
  ram[6887]  = 1;
  ram[6888]  = 1;
  ram[6889]  = 1;
  ram[6890]  = 1;
  ram[6891]  = 1;
  ram[6892]  = 1;
  ram[6893]  = 1;
  ram[6894]  = 1;
  ram[6895]  = 1;
  ram[6896]  = 1;
  ram[6897]  = 1;
  ram[6898]  = 1;
  ram[6899]  = 1;
  ram[6900]  = 1;
  ram[6901]  = 1;
  ram[6902]  = 1;
  ram[6903]  = 1;
  ram[6904]  = 1;
  ram[6905]  = 1;
  ram[6906]  = 1;
  ram[6907]  = 1;
  ram[6908]  = 1;
  ram[6909]  = 1;
  ram[6910]  = 1;
  ram[6911]  = 1;
  ram[6912]  = 1;
  ram[6913]  = 1;
  ram[6914]  = 1;
  ram[6915]  = 1;
  ram[6916]  = 1;
  ram[6917]  = 1;
  ram[6918]  = 1;
  ram[6919]  = 1;
  ram[6920]  = 1;
  ram[6921]  = 1;
  ram[6922]  = 1;
  ram[6923]  = 1;
  ram[6924]  = 1;
  ram[6925]  = 1;
  ram[6926]  = 1;
  ram[6927]  = 1;
  ram[6928]  = 1;
  ram[6929]  = 1;
  ram[6930]  = 1;
  ram[6931]  = 1;
  ram[6932]  = 1;
  ram[6933]  = 1;
  ram[6934]  = 1;
  ram[6935]  = 1;
  ram[6936]  = 1;
  ram[6937]  = 1;
  ram[6938]  = 1;
  ram[6939]  = 1;
  ram[6940]  = 1;
  ram[6941]  = 1;
  ram[6942]  = 1;
  ram[6943]  = 1;
  ram[6944]  = 1;
  ram[6945]  = 1;
  ram[6946]  = 1;
  ram[6947]  = 1;
  ram[6948]  = 1;
  ram[6949]  = 1;
  ram[6950]  = 1;
  ram[6951]  = 1;
  ram[6952]  = 1;
  ram[6953]  = 1;
  ram[6954]  = 1;
  ram[6955]  = 1;
  ram[6956]  = 1;
  ram[6957]  = 1;
  ram[6958]  = 1;
  ram[6959]  = 1;
  ram[6960]  = 1;
  ram[6961]  = 1;
  ram[6962]  = 1;
  ram[6963]  = 1;
  ram[6964]  = 1;
  ram[6965]  = 1;
  ram[6966]  = 1;
  ram[6967]  = 1;
  ram[6968]  = 1;
  ram[6969]  = 1;
  ram[6970]  = 1;
  ram[6971]  = 1;
  ram[6972]  = 1;
  ram[6973]  = 1;
  ram[6974]  = 1;
  ram[6975]  = 1;
  ram[6976]  = 1;
  ram[6977]  = 1;
  ram[6978]  = 1;
  ram[6979]  = 1;
  ram[6980]  = 1;
  ram[6981]  = 1;
  ram[6982]  = 1;
  ram[6983]  = 1;
  ram[6984]  = 1;
  ram[6985]  = 1;
  ram[6986]  = 1;
  ram[6987]  = 1;
  ram[6988]  = 1;
  ram[6989]  = 1;
  ram[6990]  = 1;
  ram[6991]  = 1;
  ram[6992]  = 1;
  ram[6993]  = 1;
  ram[6994]  = 1;
  ram[6995]  = 1;
  ram[6996]  = 1;
  ram[6997]  = 1;
  ram[6998]  = 1;
  ram[6999]  = 1;
  ram[7000]  = 0;
  ram[7001]  = 0;
  ram[7002]  = 1;
  ram[7003]  = 1;
  ram[7004]  = 1;
  ram[7005]  = 1;
  ram[7006]  = 1;
  ram[7007]  = 1;
  ram[7008]  = 1;
  ram[7009]  = 1;
  ram[7010]  = 1;
  ram[7011]  = 1;
  ram[7012]  = 1;
  ram[7013]  = 1;
  ram[7014]  = 0;
  ram[7015]  = 0;
  ram[7016]  = 0;
  ram[7017]  = 0;
  ram[7018]  = 1;
  ram[7019]  = 1;
  ram[7020]  = 1;
  ram[7021]  = 1;
  ram[7022]  = 0;
  ram[7023]  = 1;
  ram[7024]  = 1;
  ram[7025]  = 0;
  ram[7026]  = 0;
  ram[7027]  = 0;
  ram[7028]  = 1;
  ram[7029]  = 1;
  ram[7030]  = 0;
  ram[7031]  = 0;
  ram[7032]  = 0;
  ram[7033]  = 0;
  ram[7034]  = 1;
  ram[7035]  = 1;
  ram[7036]  = 1;
  ram[7037]  = 1;
  ram[7038]  = 1;
  ram[7039]  = 0;
  ram[7040]  = 0;
  ram[7041]  = 0;
  ram[7042]  = 0;
  ram[7043]  = 1;
  ram[7044]  = 1;
  ram[7045]  = 1;
  ram[7046]  = 1;
  ram[7047]  = 1;
  ram[7048]  = 1;
  ram[7049]  = 1;
  ram[7050]  = 1;
  ram[7051]  = 1;
  ram[7052]  = 0;
  ram[7053]  = 0;
  ram[7054]  = 1;
  ram[7055]  = 1;
  ram[7056]  = 1;
  ram[7057]  = 1;
  ram[7058]  = 1;
  ram[7059]  = 1;
  ram[7060]  = 1;
  ram[7061]  = 1;
  ram[7062]  = 0;
  ram[7063]  = 0;
  ram[7064]  = 1;
  ram[7065]  = 0;
  ram[7066]  = 1;
  ram[7067]  = 1;
  ram[7068]  = 1;
  ram[7069]  = 1;
  ram[7070]  = 1;
  ram[7071]  = 1;
  ram[7072]  = 0;
  ram[7073]  = 0;
  ram[7074]  = 1;
  ram[7075]  = 1;
  ram[7076]  = 1;
  ram[7077]  = 0;
  ram[7078]  = 0;
  ram[7079]  = 0;
  ram[7080]  = 0;
  ram[7081]  = 1;
  ram[7082]  = 1;
  ram[7083]  = 1;
  ram[7084]  = 1;
  ram[7085]  = 0;
  ram[7086]  = 1;
  ram[7087]  = 0;
  ram[7088]  = 0;
  ram[7089]  = 1;
  ram[7090]  = 1;
  ram[7091]  = 0;
  ram[7092]  = 0;
  ram[7093]  = 1;
  ram[7094]  = 1;
  ram[7095]  = 1;
  ram[7096]  = 1;
  ram[7097]  = 1;
  ram[7098]  = 1;
  ram[7099]  = 1;
  ram[7100]  = 1;
  ram[7101]  = 1;
  ram[7102]  = 1;
  ram[7103]  = 1;
  ram[7104]  = 1;
  ram[7105]  = 1;
  ram[7106]  = 1;
  ram[7107]  = 1;
  ram[7108]  = 1;
  ram[7109]  = 1;
  ram[7110]  = 1;
  ram[7111]  = 1;
  ram[7112]  = 1;
  ram[7113]  = 1;
  ram[7114]  = 1;
  ram[7115]  = 1;
  ram[7116]  = 1;
  ram[7117]  = 1;
  ram[7118]  = 1;
  ram[7119]  = 1;
  ram[7120]  = 1;
  ram[7121]  = 1;
  ram[7122]  = 1;
  ram[7123]  = 1;
  ram[7124]  = 1;
  ram[7125]  = 1;
  ram[7126]  = 1;
  ram[7127]  = 1;
  ram[7128]  = 1;
  ram[7129]  = 1;
  ram[7130]  = 1;
  ram[7131]  = 1;
  ram[7132]  = 1;
  ram[7133]  = 1;
  ram[7134]  = 1;
  ram[7135]  = 1;
  ram[7136]  = 1;
  ram[7137]  = 1;
  ram[7138]  = 1;
  ram[7139]  = 1;
  ram[7140]  = 1;
  ram[7141]  = 1;
  ram[7142]  = 1;
  ram[7143]  = 1;
  ram[7144]  = 1;
  ram[7145]  = 1;
  ram[7146]  = 1;
  ram[7147]  = 1;
  ram[7148]  = 1;
  ram[7149]  = 1;
  ram[7150]  = 1;
  ram[7151]  = 1;
  ram[7152]  = 1;
  ram[7153]  = 1;
  ram[7154]  = 1;
  ram[7155]  = 1;
  ram[7156]  = 1;
  ram[7157]  = 1;
  ram[7158]  = 1;
  ram[7159]  = 1;
  ram[7160]  = 1;
  ram[7161]  = 1;
  ram[7162]  = 1;
  ram[7163]  = 1;
  ram[7164]  = 1;
  ram[7165]  = 1;
  ram[7166]  = 1;
  ram[7167]  = 1;
  ram[7168]  = 1;
  ram[7169]  = 1;
  ram[7170]  = 1;
  ram[7171]  = 1;
  ram[7172]  = 1;
  ram[7173]  = 1;
  ram[7174]  = 1;
  ram[7175]  = 1;
  ram[7176]  = 1;
  ram[7177]  = 1;
  ram[7178]  = 1;
  ram[7179]  = 1;
  ram[7180]  = 1;
  ram[7181]  = 1;
  ram[7182]  = 1;
  ram[7183]  = 1;
  ram[7184]  = 1;
  ram[7185]  = 1;
  ram[7186]  = 1;
  ram[7187]  = 1;
  ram[7188]  = 1;
  ram[7189]  = 1;
  ram[7190]  = 1;
  ram[7191]  = 1;
  ram[7192]  = 1;
  ram[7193]  = 1;
  ram[7194]  = 1;
  ram[7195]  = 1;
  ram[7196]  = 1;
  ram[7197]  = 1;
  ram[7198]  = 1;
  ram[7199]  = 1;
  ram[7200]  = 1;
  ram[7201]  = 1;
  ram[7202]  = 1;
  ram[7203]  = 1;
  ram[7204]  = 1;
  ram[7205]  = 1;
  ram[7206]  = 1;
  ram[7207]  = 1;
  ram[7208]  = 1;
  ram[7209]  = 1;
  ram[7210]  = 1;
  ram[7211]  = 1;
  ram[7212]  = 1;
  ram[7213]  = 1;
  ram[7214]  = 1;
  ram[7215]  = 1;
  ram[7216]  = 1;
  ram[7217]  = 1;
  ram[7218]  = 1;
  ram[7219]  = 1;
  ram[7220]  = 1;
  ram[7221]  = 1;
  ram[7222]  = 1;
  ram[7223]  = 1;
  ram[7224]  = 1;
  ram[7225]  = 1;
  ram[7226]  = 1;
  ram[7227]  = 1;
  ram[7228]  = 1;
  ram[7229]  = 1;
  ram[7230]  = 1;
  ram[7231]  = 1;
  ram[7232]  = 1;
  ram[7233]  = 1;
  ram[7234]  = 1;
  ram[7235]  = 1;
  ram[7236]  = 1;
  ram[7237]  = 1;
  ram[7238]  = 1;
  ram[7239]  = 1;
  ram[7240]  = 1;
  ram[7241]  = 1;
  ram[7242]  = 1;
  ram[7243]  = 1;
  ram[7244]  = 1;
  ram[7245]  = 1;
  ram[7246]  = 1;
  ram[7247]  = 1;
  ram[7248]  = 1;
  ram[7249]  = 1;
  ram[7250]  = 1;
  ram[7251]  = 1;
  ram[7252]  = 1;
  ram[7253]  = 1;
  ram[7254]  = 1;
  ram[7255]  = 1;
  ram[7256]  = 1;
  ram[7257]  = 1;
  ram[7258]  = 1;
  ram[7259]  = 1;
  ram[7260]  = 1;
  ram[7261]  = 1;
  ram[7262]  = 1;
  ram[7263]  = 1;
  ram[7264]  = 1;
  ram[7265]  = 1;
  ram[7266]  = 1;
  ram[7267]  = 1;
  ram[7268]  = 1;
  ram[7269]  = 1;
  ram[7270]  = 1;
  ram[7271]  = 1;
  ram[7272]  = 1;
  ram[7273]  = 1;
  ram[7274]  = 1;
  ram[7275]  = 1;
  ram[7276]  = 1;
  ram[7277]  = 1;
  ram[7278]  = 1;
  ram[7279]  = 1;
  ram[7280]  = 1;
  ram[7281]  = 1;
  ram[7282]  = 1;
  ram[7283]  = 1;
  ram[7284]  = 1;
  ram[7285]  = 1;
  ram[7286]  = 1;
  ram[7287]  = 1;
  ram[7288]  = 1;
  ram[7289]  = 1;
  ram[7290]  = 1;
  ram[7291]  = 1;
  ram[7292]  = 1;
  ram[7293]  = 1;
  ram[7294]  = 1;
  ram[7295]  = 1;
  ram[7296]  = 1;
  ram[7297]  = 1;
  ram[7298]  = 1;
  ram[7299]  = 1;
  ram[7300]  = 0;
  ram[7301]  = 1;
  ram[7302]  = 1;
  ram[7303]  = 1;
  ram[7304]  = 1;
  ram[7305]  = 1;
  ram[7306]  = 1;
  ram[7307]  = 1;
  ram[7308]  = 1;
  ram[7309]  = 1;
  ram[7310]  = 1;
  ram[7311]  = 1;
  ram[7312]  = 1;
  ram[7313]  = 0;
  ram[7314]  = 0;
  ram[7315]  = 1;
  ram[7316]  = 1;
  ram[7317]  = 0;
  ram[7318]  = 0;
  ram[7319]  = 1;
  ram[7320]  = 1;
  ram[7321]  = 1;
  ram[7322]  = 0;
  ram[7323]  = 1;
  ram[7324]  = 0;
  ram[7325]  = 1;
  ram[7326]  = 1;
  ram[7327]  = 0;
  ram[7328]  = 0;
  ram[7329]  = 1;
  ram[7330]  = 0;
  ram[7331]  = 1;
  ram[7332]  = 0;
  ram[7333]  = 0;
  ram[7334]  = 1;
  ram[7335]  = 1;
  ram[7336]  = 1;
  ram[7337]  = 1;
  ram[7338]  = 1;
  ram[7339]  = 0;
  ram[7340]  = 1;
  ram[7341]  = 1;
  ram[7342]  = 0;
  ram[7343]  = 0;
  ram[7344]  = 1;
  ram[7345]  = 1;
  ram[7346]  = 1;
  ram[7347]  = 1;
  ram[7348]  = 1;
  ram[7349]  = 1;
  ram[7350]  = 1;
  ram[7351]  = 1;
  ram[7352]  = 0;
  ram[7353]  = 0;
  ram[7354]  = 1;
  ram[7355]  = 1;
  ram[7356]  = 1;
  ram[7357]  = 1;
  ram[7358]  = 1;
  ram[7359]  = 1;
  ram[7360]  = 1;
  ram[7361]  = 1;
  ram[7362]  = 1;
  ram[7363]  = 0;
  ram[7364]  = 1;
  ram[7365]  = 0;
  ram[7366]  = 0;
  ram[7367]  = 1;
  ram[7368]  = 1;
  ram[7369]  = 1;
  ram[7370]  = 1;
  ram[7371]  = 1;
  ram[7372]  = 0;
  ram[7373]  = 1;
  ram[7374]  = 1;
  ram[7375]  = 1;
  ram[7376]  = 0;
  ram[7377]  = 0;
  ram[7378]  = 1;
  ram[7379]  = 0;
  ram[7380]  = 0;
  ram[7381]  = 1;
  ram[7382]  = 1;
  ram[7383]  = 1;
  ram[7384]  = 1;
  ram[7385]  = 0;
  ram[7386]  = 0;
  ram[7387]  = 0;
  ram[7388]  = 1;
  ram[7389]  = 1;
  ram[7390]  = 1;
  ram[7391]  = 0;
  ram[7392]  = 0;
  ram[7393]  = 1;
  ram[7394]  = 1;
  ram[7395]  = 1;
  ram[7396]  = 1;
  ram[7397]  = 1;
  ram[7398]  = 1;
  ram[7399]  = 1;
  ram[7400]  = 1;
  ram[7401]  = 1;
  ram[7402]  = 1;
  ram[7403]  = 1;
  ram[7404]  = 1;
  ram[7405]  = 1;
  ram[7406]  = 1;
  ram[7407]  = 1;
  ram[7408]  = 1;
  ram[7409]  = 1;
  ram[7410]  = 1;
  ram[7411]  = 1;
  ram[7412]  = 1;
  ram[7413]  = 1;
  ram[7414]  = 1;
  ram[7415]  = 1;
  ram[7416]  = 1;
  ram[7417]  = 1;
  ram[7418]  = 1;
  ram[7419]  = 1;
  ram[7420]  = 1;
  ram[7421]  = 1;
  ram[7422]  = 1;
  ram[7423]  = 1;
  ram[7424]  = 1;
  ram[7425]  = 1;
  ram[7426]  = 1;
  ram[7427]  = 1;
  ram[7428]  = 1;
  ram[7429]  = 1;
  ram[7430]  = 1;
  ram[7431]  = 1;
  ram[7432]  = 1;
  ram[7433]  = 1;
  ram[7434]  = 1;
  ram[7435]  = 1;
  ram[7436]  = 1;
  ram[7437]  = 1;
  ram[7438]  = 1;
  ram[7439]  = 1;
  ram[7440]  = 1;
  ram[7441]  = 1;
  ram[7442]  = 1;
  ram[7443]  = 1;
  ram[7444]  = 1;
  ram[7445]  = 1;
  ram[7446]  = 1;
  ram[7447]  = 1;
  ram[7448]  = 1;
  ram[7449]  = 1;
  ram[7450]  = 1;
  ram[7451]  = 1;
  ram[7452]  = 1;
  ram[7453]  = 1;
  ram[7454]  = 1;
  ram[7455]  = 1;
  ram[7456]  = 1;
  ram[7457]  = 1;
  ram[7458]  = 1;
  ram[7459]  = 1;
  ram[7460]  = 1;
  ram[7461]  = 1;
  ram[7462]  = 1;
  ram[7463]  = 1;
  ram[7464]  = 1;
  ram[7465]  = 1;
  ram[7466]  = 1;
  ram[7467]  = 1;
  ram[7468]  = 1;
  ram[7469]  = 1;
  ram[7470]  = 1;
  ram[7471]  = 1;
  ram[7472]  = 1;
  ram[7473]  = 1;
  ram[7474]  = 1;
  ram[7475]  = 1;
  ram[7476]  = 1;
  ram[7477]  = 1;
  ram[7478]  = 1;
  ram[7479]  = 1;
  ram[7480]  = 1;
  ram[7481]  = 1;
  ram[7482]  = 1;
  ram[7483]  = 1;
  ram[7484]  = 1;
  ram[7485]  = 1;
  ram[7486]  = 1;
  ram[7487]  = 1;
  ram[7488]  = 1;
  ram[7489]  = 1;
  ram[7490]  = 1;
  ram[7491]  = 1;
  ram[7492]  = 1;
  ram[7493]  = 1;
  ram[7494]  = 1;
  ram[7495]  = 1;
  ram[7496]  = 1;
  ram[7497]  = 1;
  ram[7498]  = 1;
  ram[7499]  = 1;
  ram[7500]  = 1;
  ram[7501]  = 1;
  ram[7502]  = 1;
  ram[7503]  = 1;
  ram[7504]  = 1;
  ram[7505]  = 1;
  ram[7506]  = 1;
  ram[7507]  = 1;
  ram[7508]  = 1;
  ram[7509]  = 1;
  ram[7510]  = 1;
  ram[7511]  = 1;
  ram[7512]  = 1;
  ram[7513]  = 1;
  ram[7514]  = 1;
  ram[7515]  = 1;
  ram[7516]  = 1;
  ram[7517]  = 1;
  ram[7518]  = 1;
  ram[7519]  = 1;
  ram[7520]  = 1;
  ram[7521]  = 1;
  ram[7522]  = 1;
  ram[7523]  = 1;
  ram[7524]  = 1;
  ram[7525]  = 1;
  ram[7526]  = 1;
  ram[7527]  = 1;
  ram[7528]  = 1;
  ram[7529]  = 1;
  ram[7530]  = 1;
  ram[7531]  = 1;
  ram[7532]  = 1;
  ram[7533]  = 1;
  ram[7534]  = 1;
  ram[7535]  = 1;
  ram[7536]  = 1;
  ram[7537]  = 1;
  ram[7538]  = 1;
  ram[7539]  = 1;
  ram[7540]  = 1;
  ram[7541]  = 1;
  ram[7542]  = 1;
  ram[7543]  = 1;
  ram[7544]  = 1;
  ram[7545]  = 1;
  ram[7546]  = 1;
  ram[7547]  = 1;
  ram[7548]  = 1;
  ram[7549]  = 1;
  ram[7550]  = 1;
  ram[7551]  = 1;
  ram[7552]  = 1;
  ram[7553]  = 1;
  ram[7554]  = 1;
  ram[7555]  = 1;
  ram[7556]  = 1;
  ram[7557]  = 1;
  ram[7558]  = 1;
  ram[7559]  = 1;
  ram[7560]  = 1;
  ram[7561]  = 1;
  ram[7562]  = 1;
  ram[7563]  = 1;
  ram[7564]  = 1;
  ram[7565]  = 1;
  ram[7566]  = 1;
  ram[7567]  = 1;
  ram[7568]  = 1;
  ram[7569]  = 1;
  ram[7570]  = 1;
  ram[7571]  = 1;
  ram[7572]  = 1;
  ram[7573]  = 1;
  ram[7574]  = 1;
  ram[7575]  = 1;
  ram[7576]  = 1;
  ram[7577]  = 1;
  ram[7578]  = 1;
  ram[7579]  = 1;
  ram[7580]  = 1;
  ram[7581]  = 1;
  ram[7582]  = 1;
  ram[7583]  = 1;
  ram[7584]  = 1;
  ram[7585]  = 1;
  ram[7586]  = 1;
  ram[7587]  = 1;
  ram[7588]  = 1;
  ram[7589]  = 1;
  ram[7590]  = 1;
  ram[7591]  = 1;
  ram[7592]  = 1;
  ram[7593]  = 1;
  ram[7594]  = 1;
  ram[7595]  = 1;
  ram[7596]  = 1;
  ram[7597]  = 1;
  ram[7598]  = 1;
  ram[7599]  = 1;
  ram[7600]  = 0;
  ram[7601]  = 1;
  ram[7602]  = 1;
  ram[7603]  = 1;
  ram[7604]  = 1;
  ram[7605]  = 1;
  ram[7606]  = 1;
  ram[7607]  = 1;
  ram[7608]  = 1;
  ram[7609]  = 1;
  ram[7610]  = 1;
  ram[7611]  = 1;
  ram[7612]  = 1;
  ram[7613]  = 0;
  ram[7614]  = 1;
  ram[7615]  = 1;
  ram[7616]  = 1;
  ram[7617]  = 1;
  ram[7618]  = 0;
  ram[7619]  = 1;
  ram[7620]  = 1;
  ram[7621]  = 1;
  ram[7622]  = 0;
  ram[7623]  = 0;
  ram[7624]  = 1;
  ram[7625]  = 1;
  ram[7626]  = 1;
  ram[7627]  = 1;
  ram[7628]  = 0;
  ram[7629]  = 0;
  ram[7630]  = 1;
  ram[7631]  = 1;
  ram[7632]  = 1;
  ram[7633]  = 0;
  ram[7634]  = 0;
  ram[7635]  = 1;
  ram[7636]  = 1;
  ram[7637]  = 1;
  ram[7638]  = 0;
  ram[7639]  = 1;
  ram[7640]  = 1;
  ram[7641]  = 1;
  ram[7642]  = 1;
  ram[7643]  = 0;
  ram[7644]  = 0;
  ram[7645]  = 1;
  ram[7646]  = 1;
  ram[7647]  = 1;
  ram[7648]  = 1;
  ram[7649]  = 1;
  ram[7650]  = 1;
  ram[7651]  = 1;
  ram[7652]  = 0;
  ram[7653]  = 1;
  ram[7654]  = 1;
  ram[7655]  = 1;
  ram[7656]  = 1;
  ram[7657]  = 1;
  ram[7658]  = 1;
  ram[7659]  = 1;
  ram[7660]  = 1;
  ram[7661]  = 1;
  ram[7662]  = 1;
  ram[7663]  = 0;
  ram[7664]  = 1;
  ram[7665]  = 1;
  ram[7666]  = 0;
  ram[7667]  = 1;
  ram[7668]  = 1;
  ram[7669]  = 1;
  ram[7670]  = 1;
  ram[7671]  = 1;
  ram[7672]  = 0;
  ram[7673]  = 1;
  ram[7674]  = 1;
  ram[7675]  = 0;
  ram[7676]  = 0;
  ram[7677]  = 1;
  ram[7678]  = 1;
  ram[7679]  = 1;
  ram[7680]  = 0;
  ram[7681]  = 0;
  ram[7682]  = 1;
  ram[7683]  = 1;
  ram[7684]  = 1;
  ram[7685]  = 0;
  ram[7686]  = 0;
  ram[7687]  = 1;
  ram[7688]  = 1;
  ram[7689]  = 1;
  ram[7690]  = 1;
  ram[7691]  = 0;
  ram[7692]  = 0;
  ram[7693]  = 1;
  ram[7694]  = 1;
  ram[7695]  = 1;
  ram[7696]  = 1;
  ram[7697]  = 1;
  ram[7698]  = 1;
  ram[7699]  = 1;
  ram[7700]  = 1;
  ram[7701]  = 1;
  ram[7702]  = 1;
  ram[7703]  = 1;
  ram[7704]  = 1;
  ram[7705]  = 1;
  ram[7706]  = 1;
  ram[7707]  = 1;
  ram[7708]  = 1;
  ram[7709]  = 1;
  ram[7710]  = 1;
  ram[7711]  = 1;
  ram[7712]  = 1;
  ram[7713]  = 1;
  ram[7714]  = 1;
  ram[7715]  = 1;
  ram[7716]  = 1;
  ram[7717]  = 1;
  ram[7718]  = 1;
  ram[7719]  = 1;
  ram[7720]  = 1;
  ram[7721]  = 1;
  ram[7722]  = 1;
  ram[7723]  = 1;
  ram[7724]  = 1;
  ram[7725]  = 1;
  ram[7726]  = 1;
  ram[7727]  = 1;
  ram[7728]  = 1;
  ram[7729]  = 1;
  ram[7730]  = 1;
  ram[7731]  = 1;
  ram[7732]  = 1;
  ram[7733]  = 1;
  ram[7734]  = 1;
  ram[7735]  = 1;
  ram[7736]  = 1;
  ram[7737]  = 1;
  ram[7738]  = 1;
  ram[7739]  = 1;
  ram[7740]  = 1;
  ram[7741]  = 1;
  ram[7742]  = 1;
  ram[7743]  = 1;
  ram[7744]  = 1;
  ram[7745]  = 1;
  ram[7746]  = 1;
  ram[7747]  = 1;
  ram[7748]  = 1;
  ram[7749]  = 1;
  ram[7750]  = 1;
  ram[7751]  = 1;
  ram[7752]  = 1;
  ram[7753]  = 1;
  ram[7754]  = 1;
  ram[7755]  = 1;
  ram[7756]  = 1;
  ram[7757]  = 1;
  ram[7758]  = 1;
  ram[7759]  = 1;
  ram[7760]  = 1;
  ram[7761]  = 1;
  ram[7762]  = 1;
  ram[7763]  = 1;
  ram[7764]  = 1;
  ram[7765]  = 1;
  ram[7766]  = 1;
  ram[7767]  = 1;
  ram[7768]  = 1;
  ram[7769]  = 1;
  ram[7770]  = 1;
  ram[7771]  = 1;
  ram[7772]  = 1;
  ram[7773]  = 1;
  ram[7774]  = 1;
  ram[7775]  = 1;
  ram[7776]  = 1;
  ram[7777]  = 1;
  ram[7778]  = 1;
  ram[7779]  = 1;
  ram[7780]  = 1;
  ram[7781]  = 1;
  ram[7782]  = 1;
  ram[7783]  = 1;
  ram[7784]  = 1;
  ram[7785]  = 1;
  ram[7786]  = 1;
  ram[7787]  = 1;
  ram[7788]  = 1;
  ram[7789]  = 1;
  ram[7790]  = 1;
  ram[7791]  = 1;
  ram[7792]  = 1;
  ram[7793]  = 1;
  ram[7794]  = 1;
  ram[7795]  = 1;
  ram[7796]  = 1;
  ram[7797]  = 1;
  ram[7798]  = 1;
  ram[7799]  = 1;
  ram[7800]  = 1;
  ram[7801]  = 1;
  ram[7802]  = 1;
  ram[7803]  = 1;
  ram[7804]  = 1;
  ram[7805]  = 1;
  ram[7806]  = 1;
  ram[7807]  = 1;
  ram[7808]  = 1;
  ram[7809]  = 1;
  ram[7810]  = 1;
  ram[7811]  = 1;
  ram[7812]  = 1;
  ram[7813]  = 1;
  ram[7814]  = 1;
  ram[7815]  = 1;
  ram[7816]  = 1;
  ram[7817]  = 1;
  ram[7818]  = 1;
  ram[7819]  = 1;
  ram[7820]  = 1;
  ram[7821]  = 1;
  ram[7822]  = 1;
  ram[7823]  = 1;
  ram[7824]  = 1;
  ram[7825]  = 1;
  ram[7826]  = 1;
  ram[7827]  = 1;
  ram[7828]  = 1;
  ram[7829]  = 1;
  ram[7830]  = 1;
  ram[7831]  = 1;
  ram[7832]  = 1;
  ram[7833]  = 1;
  ram[7834]  = 1;
  ram[7835]  = 1;
  ram[7836]  = 1;
  ram[7837]  = 1;
  ram[7838]  = 1;
  ram[7839]  = 1;
  ram[7840]  = 1;
  ram[7841]  = 1;
  ram[7842]  = 1;
  ram[7843]  = 1;
  ram[7844]  = 1;
  ram[7845]  = 1;
  ram[7846]  = 1;
  ram[7847]  = 1;
  ram[7848]  = 1;
  ram[7849]  = 1;
  ram[7850]  = 1;
  ram[7851]  = 1;
  ram[7852]  = 1;
  ram[7853]  = 1;
  ram[7854]  = 1;
  ram[7855]  = 1;
  ram[7856]  = 1;
  ram[7857]  = 1;
  ram[7858]  = 1;
  ram[7859]  = 1;
  ram[7860]  = 1;
  ram[7861]  = 1;
  ram[7862]  = 1;
  ram[7863]  = 1;
  ram[7864]  = 1;
  ram[7865]  = 1;
  ram[7866]  = 1;
  ram[7867]  = 1;
  ram[7868]  = 1;
  ram[7869]  = 1;
  ram[7870]  = 1;
  ram[7871]  = 1;
  ram[7872]  = 1;
  ram[7873]  = 1;
  ram[7874]  = 1;
  ram[7875]  = 1;
  ram[7876]  = 1;
  ram[7877]  = 1;
  ram[7878]  = 1;
  ram[7879]  = 1;
  ram[7880]  = 1;
  ram[7881]  = 1;
  ram[7882]  = 1;
  ram[7883]  = 1;
  ram[7884]  = 1;
  ram[7885]  = 1;
  ram[7886]  = 1;
  ram[7887]  = 1;
  ram[7888]  = 1;
  ram[7889]  = 1;
  ram[7890]  = 1;
  ram[7891]  = 1;
  ram[7892]  = 1;
  ram[7893]  = 1;
  ram[7894]  = 1;
  ram[7895]  = 1;
  ram[7896]  = 1;
  ram[7897]  = 1;
  ram[7898]  = 1;
  ram[7899]  = 1;
  ram[7900]  = 0;
  ram[7901]  = 1;
  ram[7902]  = 1;
  ram[7903]  = 1;
  ram[7904]  = 1;
  ram[7905]  = 1;
  ram[7906]  = 1;
  ram[7907]  = 1;
  ram[7908]  = 1;
  ram[7909]  = 1;
  ram[7910]  = 1;
  ram[7911]  = 1;
  ram[7912]  = 1;
  ram[7913]  = 0;
  ram[7914]  = 1;
  ram[7915]  = 1;
  ram[7916]  = 1;
  ram[7917]  = 1;
  ram[7918]  = 0;
  ram[7919]  = 1;
  ram[7920]  = 1;
  ram[7921]  = 1;
  ram[7922]  = 0;
  ram[7923]  = 0;
  ram[7924]  = 1;
  ram[7925]  = 1;
  ram[7926]  = 1;
  ram[7927]  = 1;
  ram[7928]  = 0;
  ram[7929]  = 0;
  ram[7930]  = 1;
  ram[7931]  = 1;
  ram[7932]  = 1;
  ram[7933]  = 1;
  ram[7934]  = 0;
  ram[7935]  = 1;
  ram[7936]  = 1;
  ram[7937]  = 1;
  ram[7938]  = 0;
  ram[7939]  = 1;
  ram[7940]  = 1;
  ram[7941]  = 1;
  ram[7942]  = 1;
  ram[7943]  = 1;
  ram[7944]  = 0;
  ram[7945]  = 1;
  ram[7946]  = 1;
  ram[7947]  = 1;
  ram[7948]  = 1;
  ram[7949]  = 1;
  ram[7950]  = 1;
  ram[7951]  = 1;
  ram[7952]  = 0;
  ram[7953]  = 1;
  ram[7954]  = 1;
  ram[7955]  = 1;
  ram[7956]  = 1;
  ram[7957]  = 1;
  ram[7958]  = 1;
  ram[7959]  = 1;
  ram[7960]  = 1;
  ram[7961]  = 1;
  ram[7962]  = 1;
  ram[7963]  = 0;
  ram[7964]  = 1;
  ram[7965]  = 1;
  ram[7966]  = 0;
  ram[7967]  = 1;
  ram[7968]  = 1;
  ram[7969]  = 1;
  ram[7970]  = 1;
  ram[7971]  = 1;
  ram[7972]  = 0;
  ram[7973]  = 1;
  ram[7974]  = 1;
  ram[7975]  = 0;
  ram[7976]  = 1;
  ram[7977]  = 1;
  ram[7978]  = 1;
  ram[7979]  = 1;
  ram[7980]  = 1;
  ram[7981]  = 0;
  ram[7982]  = 1;
  ram[7983]  = 1;
  ram[7984]  = 1;
  ram[7985]  = 0;
  ram[7986]  = 1;
  ram[7987]  = 1;
  ram[7988]  = 1;
  ram[7989]  = 1;
  ram[7990]  = 1;
  ram[7991]  = 0;
  ram[7992]  = 0;
  ram[7993]  = 1;
  ram[7994]  = 1;
  ram[7995]  = 1;
  ram[7996]  = 1;
  ram[7997]  = 1;
  ram[7998]  = 1;
  ram[7999]  = 1;
  ram[8000]  = 1;
  ram[8001]  = 1;
  ram[8002]  = 1;
  ram[8003]  = 1;
  ram[8004]  = 1;
  ram[8005]  = 1;
  ram[8006]  = 1;
  ram[8007]  = 1;
  ram[8008]  = 1;
  ram[8009]  = 1;
  ram[8010]  = 1;
  ram[8011]  = 1;
  ram[8012]  = 1;
  ram[8013]  = 1;
  ram[8014]  = 1;
  ram[8015]  = 1;
  ram[8016]  = 1;
  ram[8017]  = 1;
  ram[8018]  = 1;
  ram[8019]  = 1;
  ram[8020]  = 1;
  ram[8021]  = 1;
  ram[8022]  = 1;
  ram[8023]  = 1;
  ram[8024]  = 1;
  ram[8025]  = 1;
  ram[8026]  = 1;
  ram[8027]  = 1;
  ram[8028]  = 1;
  ram[8029]  = 1;
  ram[8030]  = 1;
  ram[8031]  = 1;
  ram[8032]  = 1;
  ram[8033]  = 1;
  ram[8034]  = 1;
  ram[8035]  = 1;
  ram[8036]  = 1;
  ram[8037]  = 1;
  ram[8038]  = 1;
  ram[8039]  = 1;
  ram[8040]  = 1;
  ram[8041]  = 1;
  ram[8042]  = 1;
  ram[8043]  = 1;
  ram[8044]  = 1;
  ram[8045]  = 1;
  ram[8046]  = 1;
  ram[8047]  = 1;
  ram[8048]  = 1;
  ram[8049]  = 1;
  ram[8050]  = 1;
  ram[8051]  = 1;
  ram[8052]  = 1;
  ram[8053]  = 1;
  ram[8054]  = 1;
  ram[8055]  = 1;
  ram[8056]  = 1;
  ram[8057]  = 1;
  ram[8058]  = 1;
  ram[8059]  = 1;
  ram[8060]  = 1;
  ram[8061]  = 1;
  ram[8062]  = 1;
  ram[8063]  = 1;
  ram[8064]  = 1;
  ram[8065]  = 1;
  ram[8066]  = 1;
  ram[8067]  = 1;
  ram[8068]  = 1;
  ram[8069]  = 1;
  ram[8070]  = 1;
  ram[8071]  = 1;
  ram[8072]  = 1;
  ram[8073]  = 1;
  ram[8074]  = 1;
  ram[8075]  = 1;
  ram[8076]  = 1;
  ram[8077]  = 1;
  ram[8078]  = 1;
  ram[8079]  = 1;
  ram[8080]  = 1;
  ram[8081]  = 1;
  ram[8082]  = 1;
  ram[8083]  = 1;
  ram[8084]  = 1;
  ram[8085]  = 1;
  ram[8086]  = 1;
  ram[8087]  = 1;
  ram[8088]  = 1;
  ram[8089]  = 1;
  ram[8090]  = 1;
  ram[8091]  = 1;
  ram[8092]  = 1;
  ram[8093]  = 1;
  ram[8094]  = 1;
  ram[8095]  = 1;
  ram[8096]  = 1;
  ram[8097]  = 1;
  ram[8098]  = 1;
  ram[8099]  = 1;
  ram[8100]  = 1;
  ram[8101]  = 1;
  ram[8102]  = 1;
  ram[8103]  = 1;
  ram[8104]  = 1;
  ram[8105]  = 1;
  ram[8106]  = 1;
  ram[8107]  = 1;
  ram[8108]  = 1;
  ram[8109]  = 1;
  ram[8110]  = 1;
  ram[8111]  = 1;
  ram[8112]  = 1;
  ram[8113]  = 1;
  ram[8114]  = 1;
  ram[8115]  = 1;
  ram[8116]  = 1;
  ram[8117]  = 1;
  ram[8118]  = 1;
  ram[8119]  = 1;
  ram[8120]  = 1;
  ram[8121]  = 1;
  ram[8122]  = 1;
  ram[8123]  = 1;
  ram[8124]  = 1;
  ram[8125]  = 1;
  ram[8126]  = 1;
  ram[8127]  = 1;
  ram[8128]  = 1;
  ram[8129]  = 1;
  ram[8130]  = 1;
  ram[8131]  = 1;
  ram[8132]  = 1;
  ram[8133]  = 1;
  ram[8134]  = 1;
  ram[8135]  = 1;
  ram[8136]  = 1;
  ram[8137]  = 1;
  ram[8138]  = 1;
  ram[8139]  = 1;
  ram[8140]  = 1;
  ram[8141]  = 1;
  ram[8142]  = 1;
  ram[8143]  = 1;
  ram[8144]  = 1;
  ram[8145]  = 1;
  ram[8146]  = 1;
  ram[8147]  = 1;
  ram[8148]  = 1;
  ram[8149]  = 1;
  ram[8150]  = 1;
  ram[8151]  = 1;
  ram[8152]  = 1;
  ram[8153]  = 1;
  ram[8154]  = 1;
  ram[8155]  = 1;
  ram[8156]  = 1;
  ram[8157]  = 1;
  ram[8158]  = 1;
  ram[8159]  = 1;
  ram[8160]  = 1;
  ram[8161]  = 1;
  ram[8162]  = 1;
  ram[8163]  = 1;
  ram[8164]  = 1;
  ram[8165]  = 1;
  ram[8166]  = 1;
  ram[8167]  = 1;
  ram[8168]  = 1;
  ram[8169]  = 1;
  ram[8170]  = 1;
  ram[8171]  = 1;
  ram[8172]  = 1;
  ram[8173]  = 1;
  ram[8174]  = 1;
  ram[8175]  = 1;
  ram[8176]  = 1;
  ram[8177]  = 1;
  ram[8178]  = 1;
  ram[8179]  = 1;
  ram[8180]  = 1;
  ram[8181]  = 1;
  ram[8182]  = 1;
  ram[8183]  = 1;
  ram[8184]  = 1;
  ram[8185]  = 1;
  ram[8186]  = 1;
  ram[8187]  = 1;
  ram[8188]  = 1;
  ram[8189]  = 1;
  ram[8190]  = 1;
  ram[8191]  = 1;
  ram[8192]  = 1;
  ram[8193]  = 1;
  ram[8194]  = 1;
  ram[8195]  = 1;
  ram[8196]  = 1;
  ram[8197]  = 1;
  ram[8198]  = 1;
  ram[8199]  = 1;
  ram[8200]  = 0;
  ram[8201]  = 1;
  ram[8202]  = 1;
  ram[8203]  = 1;
  ram[8204]  = 1;
  ram[8205]  = 1;
  ram[8206]  = 1;
  ram[8207]  = 1;
  ram[8208]  = 1;
  ram[8209]  = 1;
  ram[8210]  = 1;
  ram[8211]  = 1;
  ram[8212]  = 1;
  ram[8213]  = 1;
  ram[8214]  = 1;
  ram[8215]  = 1;
  ram[8216]  = 1;
  ram[8217]  = 1;
  ram[8218]  = 0;
  ram[8219]  = 1;
  ram[8220]  = 1;
  ram[8221]  = 1;
  ram[8222]  = 0;
  ram[8223]  = 0;
  ram[8224]  = 1;
  ram[8225]  = 1;
  ram[8226]  = 1;
  ram[8227]  = 1;
  ram[8228]  = 0;
  ram[8229]  = 1;
  ram[8230]  = 1;
  ram[8231]  = 1;
  ram[8232]  = 1;
  ram[8233]  = 1;
  ram[8234]  = 0;
  ram[8235]  = 1;
  ram[8236]  = 1;
  ram[8237]  = 1;
  ram[8238]  = 0;
  ram[8239]  = 1;
  ram[8240]  = 1;
  ram[8241]  = 1;
  ram[8242]  = 1;
  ram[8243]  = 1;
  ram[8244]  = 0;
  ram[8245]  = 1;
  ram[8246]  = 1;
  ram[8247]  = 1;
  ram[8248]  = 1;
  ram[8249]  = 1;
  ram[8250]  = 1;
  ram[8251]  = 1;
  ram[8252]  = 0;
  ram[8253]  = 1;
  ram[8254]  = 1;
  ram[8255]  = 1;
  ram[8256]  = 1;
  ram[8257]  = 1;
  ram[8258]  = 1;
  ram[8259]  = 1;
  ram[8260]  = 1;
  ram[8261]  = 1;
  ram[8262]  = 1;
  ram[8263]  = 0;
  ram[8264]  = 1;
  ram[8265]  = 1;
  ram[8266]  = 0;
  ram[8267]  = 1;
  ram[8268]  = 1;
  ram[8269]  = 1;
  ram[8270]  = 1;
  ram[8271]  = 0;
  ram[8272]  = 0;
  ram[8273]  = 1;
  ram[8274]  = 1;
  ram[8275]  = 0;
  ram[8276]  = 1;
  ram[8277]  = 1;
  ram[8278]  = 1;
  ram[8279]  = 1;
  ram[8280]  = 1;
  ram[8281]  = 0;
  ram[8282]  = 1;
  ram[8283]  = 1;
  ram[8284]  = 1;
  ram[8285]  = 0;
  ram[8286]  = 1;
  ram[8287]  = 1;
  ram[8288]  = 1;
  ram[8289]  = 1;
  ram[8290]  = 1;
  ram[8291]  = 1;
  ram[8292]  = 0;
  ram[8293]  = 1;
  ram[8294]  = 1;
  ram[8295]  = 1;
  ram[8296]  = 1;
  ram[8297]  = 1;
  ram[8298]  = 1;
  ram[8299]  = 1;
  ram[8300]  = 1;
  ram[8301]  = 1;
  ram[8302]  = 1;
  ram[8303]  = 1;
  ram[8304]  = 1;
  ram[8305]  = 1;
  ram[8306]  = 1;
  ram[8307]  = 1;
  ram[8308]  = 1;
  ram[8309]  = 1;
  ram[8310]  = 1;
  ram[8311]  = 1;
  ram[8312]  = 1;
  ram[8313]  = 1;
  ram[8314]  = 1;
  ram[8315]  = 1;
  ram[8316]  = 1;
  ram[8317]  = 1;
  ram[8318]  = 1;
  ram[8319]  = 1;
  ram[8320]  = 1;
  ram[8321]  = 1;
  ram[8322]  = 1;
  ram[8323]  = 1;
  ram[8324]  = 1;
  ram[8325]  = 1;
  ram[8326]  = 1;
  ram[8327]  = 1;
  ram[8328]  = 1;
  ram[8329]  = 1;
  ram[8330]  = 1;
  ram[8331]  = 1;
  ram[8332]  = 1;
  ram[8333]  = 1;
  ram[8334]  = 1;
  ram[8335]  = 1;
  ram[8336]  = 1;
  ram[8337]  = 1;
  ram[8338]  = 1;
  ram[8339]  = 1;
  ram[8340]  = 1;
  ram[8341]  = 1;
  ram[8342]  = 1;
  ram[8343]  = 1;
  ram[8344]  = 1;
  ram[8345]  = 1;
  ram[8346]  = 1;
  ram[8347]  = 1;
  ram[8348]  = 1;
  ram[8349]  = 1;
  ram[8350]  = 1;
  ram[8351]  = 1;
  ram[8352]  = 1;
  ram[8353]  = 1;
  ram[8354]  = 1;
  ram[8355]  = 1;
  ram[8356]  = 1;
  ram[8357]  = 1;
  ram[8358]  = 1;
  ram[8359]  = 1;
  ram[8360]  = 1;
  ram[8361]  = 1;
  ram[8362]  = 1;
  ram[8363]  = 1;
  ram[8364]  = 1;
  ram[8365]  = 1;
  ram[8366]  = 1;
  ram[8367]  = 1;
  ram[8368]  = 1;
  ram[8369]  = 1;
  ram[8370]  = 1;
  ram[8371]  = 1;
  ram[8372]  = 1;
  ram[8373]  = 1;
  ram[8374]  = 1;
  ram[8375]  = 1;
  ram[8376]  = 1;
  ram[8377]  = 1;
  ram[8378]  = 1;
  ram[8379]  = 1;
  ram[8380]  = 1;
  ram[8381]  = 1;
  ram[8382]  = 1;
  ram[8383]  = 1;
  ram[8384]  = 1;
  ram[8385]  = 1;
  ram[8386]  = 1;
  ram[8387]  = 1;
  ram[8388]  = 1;
  ram[8389]  = 1;
  ram[8390]  = 1;
  ram[8391]  = 1;
  ram[8392]  = 1;
  ram[8393]  = 1;
  ram[8394]  = 1;
  ram[8395]  = 1;
  ram[8396]  = 1;
  ram[8397]  = 1;
  ram[8398]  = 1;
  ram[8399]  = 1;
  ram[8400]  = 1;
  ram[8401]  = 1;
  ram[8402]  = 1;
  ram[8403]  = 1;
  ram[8404]  = 1;
  ram[8405]  = 1;
  ram[8406]  = 1;
  ram[8407]  = 1;
  ram[8408]  = 1;
  ram[8409]  = 1;
  ram[8410]  = 1;
  ram[8411]  = 1;
  ram[8412]  = 1;
  ram[8413]  = 1;
  ram[8414]  = 1;
  ram[8415]  = 1;
  ram[8416]  = 1;
  ram[8417]  = 1;
  ram[8418]  = 1;
  ram[8419]  = 1;
  ram[8420]  = 1;
  ram[8421]  = 1;
  ram[8422]  = 1;
  ram[8423]  = 1;
  ram[8424]  = 1;
  ram[8425]  = 1;
  ram[8426]  = 1;
  ram[8427]  = 1;
  ram[8428]  = 1;
  ram[8429]  = 1;
  ram[8430]  = 1;
  ram[8431]  = 1;
  ram[8432]  = 1;
  ram[8433]  = 1;
  ram[8434]  = 1;
  ram[8435]  = 1;
  ram[8436]  = 1;
  ram[8437]  = 1;
  ram[8438]  = 1;
  ram[8439]  = 1;
  ram[8440]  = 1;
  ram[8441]  = 1;
  ram[8442]  = 1;
  ram[8443]  = 1;
  ram[8444]  = 1;
  ram[8445]  = 1;
  ram[8446]  = 1;
  ram[8447]  = 1;
  ram[8448]  = 1;
  ram[8449]  = 1;
  ram[8450]  = 1;
  ram[8451]  = 1;
  ram[8452]  = 1;
  ram[8453]  = 1;
  ram[8454]  = 1;
  ram[8455]  = 1;
  ram[8456]  = 1;
  ram[8457]  = 1;
  ram[8458]  = 1;
  ram[8459]  = 1;
  ram[8460]  = 1;
  ram[8461]  = 1;
  ram[8462]  = 1;
  ram[8463]  = 1;
  ram[8464]  = 1;
  ram[8465]  = 1;
  ram[8466]  = 1;
  ram[8467]  = 1;
  ram[8468]  = 1;
  ram[8469]  = 1;
  ram[8470]  = 1;
  ram[8471]  = 1;
  ram[8472]  = 1;
  ram[8473]  = 1;
  ram[8474]  = 1;
  ram[8475]  = 1;
  ram[8476]  = 1;
  ram[8477]  = 1;
  ram[8478]  = 1;
  ram[8479]  = 1;
  ram[8480]  = 1;
  ram[8481]  = 1;
  ram[8482]  = 1;
  ram[8483]  = 1;
  ram[8484]  = 1;
  ram[8485]  = 1;
  ram[8486]  = 1;
  ram[8487]  = 1;
  ram[8488]  = 1;
  ram[8489]  = 1;
  ram[8490]  = 1;
  ram[8491]  = 1;
  ram[8492]  = 1;
  ram[8493]  = 1;
  ram[8494]  = 1;
  ram[8495]  = 1;
  ram[8496]  = 1;
  ram[8497]  = 1;
  ram[8498]  = 1;
  ram[8499]  = 1;
  ram[8500]  = 0;
  ram[8501]  = 1;
  ram[8502]  = 1;
  ram[8503]  = 1;
  ram[8504]  = 1;
  ram[8505]  = 1;
  ram[8506]  = 0;
  ram[8507]  = 0;
  ram[8508]  = 0;
  ram[8509]  = 0;
  ram[8510]  = 1;
  ram[8511]  = 1;
  ram[8512]  = 1;
  ram[8513]  = 1;
  ram[8514]  = 1;
  ram[8515]  = 1;
  ram[8516]  = 1;
  ram[8517]  = 1;
  ram[8518]  = 0;
  ram[8519]  = 1;
  ram[8520]  = 1;
  ram[8521]  = 1;
  ram[8522]  = 0;
  ram[8523]  = 0;
  ram[8524]  = 1;
  ram[8525]  = 1;
  ram[8526]  = 1;
  ram[8527]  = 1;
  ram[8528]  = 0;
  ram[8529]  = 1;
  ram[8530]  = 1;
  ram[8531]  = 1;
  ram[8532]  = 1;
  ram[8533]  = 1;
  ram[8534]  = 0;
  ram[8535]  = 1;
  ram[8536]  = 1;
  ram[8537]  = 0;
  ram[8538]  = 0;
  ram[8539]  = 1;
  ram[8540]  = 1;
  ram[8541]  = 1;
  ram[8542]  = 1;
  ram[8543]  = 1;
  ram[8544]  = 0;
  ram[8545]  = 1;
  ram[8546]  = 1;
  ram[8547]  = 1;
  ram[8548]  = 1;
  ram[8549]  = 1;
  ram[8550]  = 1;
  ram[8551]  = 1;
  ram[8552]  = 0;
  ram[8553]  = 1;
  ram[8554]  = 1;
  ram[8555]  = 1;
  ram[8556]  = 1;
  ram[8557]  = 1;
  ram[8558]  = 1;
  ram[8559]  = 1;
  ram[8560]  = 1;
  ram[8561]  = 1;
  ram[8562]  = 1;
  ram[8563]  = 0;
  ram[8564]  = 1;
  ram[8565]  = 1;
  ram[8566]  = 0;
  ram[8567]  = 0;
  ram[8568]  = 1;
  ram[8569]  = 1;
  ram[8570]  = 1;
  ram[8571]  = 0;
  ram[8572]  = 1;
  ram[8573]  = 1;
  ram[8574]  = 1;
  ram[8575]  = 0;
  ram[8576]  = 1;
  ram[8577]  = 1;
  ram[8578]  = 1;
  ram[8579]  = 1;
  ram[8580]  = 1;
  ram[8581]  = 0;
  ram[8582]  = 1;
  ram[8583]  = 1;
  ram[8584]  = 1;
  ram[8585]  = 0;
  ram[8586]  = 1;
  ram[8587]  = 1;
  ram[8588]  = 1;
  ram[8589]  = 1;
  ram[8590]  = 1;
  ram[8591]  = 1;
  ram[8592]  = 0;
  ram[8593]  = 1;
  ram[8594]  = 1;
  ram[8595]  = 1;
  ram[8596]  = 1;
  ram[8597]  = 1;
  ram[8598]  = 1;
  ram[8599]  = 1;
  ram[8600]  = 1;
  ram[8601]  = 1;
  ram[8602]  = 1;
  ram[8603]  = 1;
  ram[8604]  = 1;
  ram[8605]  = 1;
  ram[8606]  = 1;
  ram[8607]  = 1;
  ram[8608]  = 1;
  ram[8609]  = 1;
  ram[8610]  = 1;
  ram[8611]  = 1;
  ram[8612]  = 1;
  ram[8613]  = 1;
  ram[8614]  = 1;
  ram[8615]  = 1;
  ram[8616]  = 1;
  ram[8617]  = 1;
  ram[8618]  = 1;
  ram[8619]  = 1;
  ram[8620]  = 1;
  ram[8621]  = 1;
  ram[8622]  = 1;
  ram[8623]  = 1;
  ram[8624]  = 1;
  ram[8625]  = 1;
  ram[8626]  = 1;
  ram[8627]  = 1;
  ram[8628]  = 1;
  ram[8629]  = 1;
  ram[8630]  = 1;
  ram[8631]  = 1;
  ram[8632]  = 1;
  ram[8633]  = 1;
  ram[8634]  = 1;
  ram[8635]  = 1;
  ram[8636]  = 1;
  ram[8637]  = 1;
  ram[8638]  = 1;
  ram[8639]  = 1;
  ram[8640]  = 1;
  ram[8641]  = 1;
  ram[8642]  = 1;
  ram[8643]  = 1;
  ram[8644]  = 1;
  ram[8645]  = 1;
  ram[8646]  = 1;
  ram[8647]  = 1;
  ram[8648]  = 1;
  ram[8649]  = 1;
  ram[8650]  = 1;
  ram[8651]  = 1;
  ram[8652]  = 1;
  ram[8653]  = 1;
  ram[8654]  = 1;
  ram[8655]  = 1;
  ram[8656]  = 1;
  ram[8657]  = 1;
  ram[8658]  = 1;
  ram[8659]  = 1;
  ram[8660]  = 1;
  ram[8661]  = 1;
  ram[8662]  = 1;
  ram[8663]  = 1;
  ram[8664]  = 1;
  ram[8665]  = 1;
  ram[8666]  = 1;
  ram[8667]  = 1;
  ram[8668]  = 1;
  ram[8669]  = 1;
  ram[8670]  = 1;
  ram[8671]  = 1;
  ram[8672]  = 1;
  ram[8673]  = 1;
  ram[8674]  = 1;
  ram[8675]  = 1;
  ram[8676]  = 1;
  ram[8677]  = 1;
  ram[8678]  = 1;
  ram[8679]  = 1;
  ram[8680]  = 1;
  ram[8681]  = 1;
  ram[8682]  = 1;
  ram[8683]  = 1;
  ram[8684]  = 1;
  ram[8685]  = 1;
  ram[8686]  = 1;
  ram[8687]  = 1;
  ram[8688]  = 1;
  ram[8689]  = 1;
  ram[8690]  = 1;
  ram[8691]  = 1;
  ram[8692]  = 1;
  ram[8693]  = 1;
  ram[8694]  = 1;
  ram[8695]  = 1;
  ram[8696]  = 1;
  ram[8697]  = 1;
  ram[8698]  = 1;
  ram[8699]  = 1;
  ram[8700]  = 1;
  ram[8701]  = 1;
  ram[8702]  = 1;
  ram[8703]  = 1;
  ram[8704]  = 1;
  ram[8705]  = 1;
  ram[8706]  = 1;
  ram[8707]  = 1;
  ram[8708]  = 1;
  ram[8709]  = 1;
  ram[8710]  = 1;
  ram[8711]  = 1;
  ram[8712]  = 1;
  ram[8713]  = 1;
  ram[8714]  = 1;
  ram[8715]  = 1;
  ram[8716]  = 1;
  ram[8717]  = 1;
  ram[8718]  = 1;
  ram[8719]  = 1;
  ram[8720]  = 1;
  ram[8721]  = 1;
  ram[8722]  = 1;
  ram[8723]  = 1;
  ram[8724]  = 1;
  ram[8725]  = 1;
  ram[8726]  = 1;
  ram[8727]  = 1;
  ram[8728]  = 1;
  ram[8729]  = 1;
  ram[8730]  = 1;
  ram[8731]  = 1;
  ram[8732]  = 1;
  ram[8733]  = 1;
  ram[8734]  = 1;
  ram[8735]  = 1;
  ram[8736]  = 1;
  ram[8737]  = 1;
  ram[8738]  = 1;
  ram[8739]  = 1;
  ram[8740]  = 1;
  ram[8741]  = 1;
  ram[8742]  = 1;
  ram[8743]  = 1;
  ram[8744]  = 1;
  ram[8745]  = 1;
  ram[8746]  = 1;
  ram[8747]  = 1;
  ram[8748]  = 1;
  ram[8749]  = 1;
  ram[8750]  = 1;
  ram[8751]  = 1;
  ram[8752]  = 1;
  ram[8753]  = 1;
  ram[8754]  = 1;
  ram[8755]  = 1;
  ram[8756]  = 1;
  ram[8757]  = 1;
  ram[8758]  = 1;
  ram[8759]  = 1;
  ram[8760]  = 1;
  ram[8761]  = 1;
  ram[8762]  = 1;
  ram[8763]  = 1;
  ram[8764]  = 1;
  ram[8765]  = 1;
  ram[8766]  = 1;
  ram[8767]  = 1;
  ram[8768]  = 1;
  ram[8769]  = 1;
  ram[8770]  = 1;
  ram[8771]  = 1;
  ram[8772]  = 1;
  ram[8773]  = 1;
  ram[8774]  = 1;
  ram[8775]  = 1;
  ram[8776]  = 1;
  ram[8777]  = 1;
  ram[8778]  = 1;
  ram[8779]  = 1;
  ram[8780]  = 1;
  ram[8781]  = 1;
  ram[8782]  = 1;
  ram[8783]  = 1;
  ram[8784]  = 1;
  ram[8785]  = 1;
  ram[8786]  = 1;
  ram[8787]  = 1;
  ram[8788]  = 1;
  ram[8789]  = 1;
  ram[8790]  = 1;
  ram[8791]  = 1;
  ram[8792]  = 1;
  ram[8793]  = 1;
  ram[8794]  = 1;
  ram[8795]  = 1;
  ram[8796]  = 1;
  ram[8797]  = 1;
  ram[8798]  = 1;
  ram[8799]  = 1;
  ram[8800]  = 0;
  ram[8801]  = 1;
  ram[8802]  = 1;
  ram[8803]  = 1;
  ram[8804]  = 1;
  ram[8805]  = 1;
  ram[8806]  = 0;
  ram[8807]  = 0;
  ram[8808]  = 0;
  ram[8809]  = 0;
  ram[8810]  = 1;
  ram[8811]  = 1;
  ram[8812]  = 1;
  ram[8813]  = 1;
  ram[8814]  = 1;
  ram[8815]  = 1;
  ram[8816]  = 0;
  ram[8817]  = 0;
  ram[8818]  = 0;
  ram[8819]  = 1;
  ram[8820]  = 1;
  ram[8821]  = 1;
  ram[8822]  = 0;
  ram[8823]  = 0;
  ram[8824]  = 1;
  ram[8825]  = 1;
  ram[8826]  = 1;
  ram[8827]  = 1;
  ram[8828]  = 0;
  ram[8829]  = 1;
  ram[8830]  = 1;
  ram[8831]  = 1;
  ram[8832]  = 1;
  ram[8833]  = 1;
  ram[8834]  = 0;
  ram[8835]  = 1;
  ram[8836]  = 1;
  ram[8837]  = 0;
  ram[8838]  = 0;
  ram[8839]  = 1;
  ram[8840]  = 1;
  ram[8841]  = 1;
  ram[8842]  = 1;
  ram[8843]  = 1;
  ram[8844]  = 0;
  ram[8845]  = 1;
  ram[8846]  = 1;
  ram[8847]  = 1;
  ram[8848]  = 1;
  ram[8849]  = 1;
  ram[8850]  = 1;
  ram[8851]  = 1;
  ram[8852]  = 0;
  ram[8853]  = 1;
  ram[8854]  = 1;
  ram[8855]  = 1;
  ram[8856]  = 1;
  ram[8857]  = 1;
  ram[8858]  = 1;
  ram[8859]  = 1;
  ram[8860]  = 1;
  ram[8861]  = 1;
  ram[8862]  = 1;
  ram[8863]  = 0;
  ram[8864]  = 1;
  ram[8865]  = 1;
  ram[8866]  = 0;
  ram[8867]  = 0;
  ram[8868]  = 1;
  ram[8869]  = 1;
  ram[8870]  = 1;
  ram[8871]  = 0;
  ram[8872]  = 1;
  ram[8873]  = 1;
  ram[8874]  = 1;
  ram[8875]  = 0;
  ram[8876]  = 1;
  ram[8877]  = 1;
  ram[8878]  = 1;
  ram[8879]  = 1;
  ram[8880]  = 1;
  ram[8881]  = 0;
  ram[8882]  = 0;
  ram[8883]  = 1;
  ram[8884]  = 1;
  ram[8885]  = 0;
  ram[8886]  = 1;
  ram[8887]  = 1;
  ram[8888]  = 1;
  ram[8889]  = 1;
  ram[8890]  = 1;
  ram[8891]  = 1;
  ram[8892]  = 0;
  ram[8893]  = 1;
  ram[8894]  = 1;
  ram[8895]  = 1;
  ram[8896]  = 1;
  ram[8897]  = 1;
  ram[8898]  = 1;
  ram[8899]  = 1;
  ram[8900]  = 1;
  ram[8901]  = 1;
  ram[8902]  = 1;
  ram[8903]  = 1;
  ram[8904]  = 1;
  ram[8905]  = 1;
  ram[8906]  = 1;
  ram[8907]  = 1;
  ram[8908]  = 1;
  ram[8909]  = 1;
  ram[8910]  = 1;
  ram[8911]  = 1;
  ram[8912]  = 1;
  ram[8913]  = 1;
  ram[8914]  = 1;
  ram[8915]  = 1;
  ram[8916]  = 1;
  ram[8917]  = 1;
  ram[8918]  = 1;
  ram[8919]  = 1;
  ram[8920]  = 1;
  ram[8921]  = 1;
  ram[8922]  = 1;
  ram[8923]  = 1;
  ram[8924]  = 1;
  ram[8925]  = 1;
  ram[8926]  = 1;
  ram[8927]  = 1;
  ram[8928]  = 1;
  ram[8929]  = 1;
  ram[8930]  = 1;
  ram[8931]  = 1;
  ram[8932]  = 1;
  ram[8933]  = 1;
  ram[8934]  = 1;
  ram[8935]  = 1;
  ram[8936]  = 1;
  ram[8937]  = 1;
  ram[8938]  = 1;
  ram[8939]  = 1;
  ram[8940]  = 1;
  ram[8941]  = 1;
  ram[8942]  = 1;
  ram[8943]  = 1;
  ram[8944]  = 1;
  ram[8945]  = 1;
  ram[8946]  = 1;
  ram[8947]  = 1;
  ram[8948]  = 1;
  ram[8949]  = 1;
  ram[8950]  = 1;
  ram[8951]  = 1;
  ram[8952]  = 1;
  ram[8953]  = 1;
  ram[8954]  = 1;
  ram[8955]  = 1;
  ram[8956]  = 1;
  ram[8957]  = 1;
  ram[8958]  = 1;
  ram[8959]  = 1;
  ram[8960]  = 1;
  ram[8961]  = 1;
  ram[8962]  = 1;
  ram[8963]  = 1;
  ram[8964]  = 1;
  ram[8965]  = 1;
  ram[8966]  = 1;
  ram[8967]  = 1;
  ram[8968]  = 1;
  ram[8969]  = 1;
  ram[8970]  = 1;
  ram[8971]  = 1;
  ram[8972]  = 1;
  ram[8973]  = 1;
  ram[8974]  = 1;
  ram[8975]  = 1;
  ram[8976]  = 1;
  ram[8977]  = 1;
  ram[8978]  = 1;
  ram[8979]  = 1;
  ram[8980]  = 1;
  ram[8981]  = 1;
  ram[8982]  = 1;
  ram[8983]  = 1;
  ram[8984]  = 1;
  ram[8985]  = 1;
  ram[8986]  = 1;
  ram[8987]  = 1;
  ram[8988]  = 1;
  ram[8989]  = 1;
  ram[8990]  = 1;
  ram[8991]  = 1;
  ram[8992]  = 1;
  ram[8993]  = 1;
  ram[8994]  = 1;
  ram[8995]  = 1;
  ram[8996]  = 1;
  ram[8997]  = 1;
  ram[8998]  = 1;
  ram[8999]  = 1;
  ram[9000]  = 1;
  ram[9001]  = 1;
  ram[9002]  = 1;
  ram[9003]  = 1;
  ram[9004]  = 1;
  ram[9005]  = 1;
  ram[9006]  = 1;
  ram[9007]  = 1;
  ram[9008]  = 1;
  ram[9009]  = 1;
  ram[9010]  = 1;
  ram[9011]  = 1;
  ram[9012]  = 1;
  ram[9013]  = 1;
  ram[9014]  = 1;
  ram[9015]  = 1;
  ram[9016]  = 1;
  ram[9017]  = 1;
  ram[9018]  = 1;
  ram[9019]  = 1;
  ram[9020]  = 1;
  ram[9021]  = 1;
  ram[9022]  = 1;
  ram[9023]  = 1;
  ram[9024]  = 1;
  ram[9025]  = 1;
  ram[9026]  = 1;
  ram[9027]  = 1;
  ram[9028]  = 1;
  ram[9029]  = 1;
  ram[9030]  = 1;
  ram[9031]  = 1;
  ram[9032]  = 1;
  ram[9033]  = 1;
  ram[9034]  = 1;
  ram[9035]  = 1;
  ram[9036]  = 1;
  ram[9037]  = 1;
  ram[9038]  = 1;
  ram[9039]  = 1;
  ram[9040]  = 1;
  ram[9041]  = 1;
  ram[9042]  = 1;
  ram[9043]  = 1;
  ram[9044]  = 1;
  ram[9045]  = 1;
  ram[9046]  = 1;
  ram[9047]  = 1;
  ram[9048]  = 1;
  ram[9049]  = 1;
  ram[9050]  = 1;
  ram[9051]  = 1;
  ram[9052]  = 1;
  ram[9053]  = 1;
  ram[9054]  = 1;
  ram[9055]  = 1;
  ram[9056]  = 1;
  ram[9057]  = 1;
  ram[9058]  = 1;
  ram[9059]  = 1;
  ram[9060]  = 1;
  ram[9061]  = 1;
  ram[9062]  = 1;
  ram[9063]  = 1;
  ram[9064]  = 1;
  ram[9065]  = 1;
  ram[9066]  = 1;
  ram[9067]  = 1;
  ram[9068]  = 1;
  ram[9069]  = 1;
  ram[9070]  = 1;
  ram[9071]  = 1;
  ram[9072]  = 1;
  ram[9073]  = 1;
  ram[9074]  = 1;
  ram[9075]  = 1;
  ram[9076]  = 1;
  ram[9077]  = 1;
  ram[9078]  = 1;
  ram[9079]  = 1;
  ram[9080]  = 1;
  ram[9081]  = 1;
  ram[9082]  = 1;
  ram[9083]  = 1;
  ram[9084]  = 1;
  ram[9085]  = 1;
  ram[9086]  = 1;
  ram[9087]  = 1;
  ram[9088]  = 1;
  ram[9089]  = 1;
  ram[9090]  = 1;
  ram[9091]  = 1;
  ram[9092]  = 1;
  ram[9093]  = 1;
  ram[9094]  = 1;
  ram[9095]  = 1;
  ram[9096]  = 1;
  ram[9097]  = 1;
  ram[9098]  = 1;
  ram[9099]  = 1;
  ram[9100]  = 0;
  ram[9101]  = 1;
  ram[9102]  = 1;
  ram[9103]  = 1;
  ram[9104]  = 1;
  ram[9105]  = 1;
  ram[9106]  = 1;
  ram[9107]  = 1;
  ram[9108]  = 1;
  ram[9109]  = 0;
  ram[9110]  = 1;
  ram[9111]  = 1;
  ram[9112]  = 1;
  ram[9113]  = 1;
  ram[9114]  = 0;
  ram[9115]  = 0;
  ram[9116]  = 0;
  ram[9117]  = 0;
  ram[9118]  = 0;
  ram[9119]  = 1;
  ram[9120]  = 1;
  ram[9121]  = 1;
  ram[9122]  = 0;
  ram[9123]  = 0;
  ram[9124]  = 1;
  ram[9125]  = 1;
  ram[9126]  = 1;
  ram[9127]  = 1;
  ram[9128]  = 0;
  ram[9129]  = 1;
  ram[9130]  = 1;
  ram[9131]  = 1;
  ram[9132]  = 1;
  ram[9133]  = 1;
  ram[9134]  = 0;
  ram[9135]  = 1;
  ram[9136]  = 1;
  ram[9137]  = 0;
  ram[9138]  = 0;
  ram[9139]  = 0;
  ram[9140]  = 0;
  ram[9141]  = 0;
  ram[9142]  = 0;
  ram[9143]  = 0;
  ram[9144]  = 0;
  ram[9145]  = 1;
  ram[9146]  = 1;
  ram[9147]  = 1;
  ram[9148]  = 1;
  ram[9149]  = 1;
  ram[9150]  = 1;
  ram[9151]  = 1;
  ram[9152]  = 0;
  ram[9153]  = 1;
  ram[9154]  = 1;
  ram[9155]  = 1;
  ram[9156]  = 1;
  ram[9157]  = 1;
  ram[9158]  = 1;
  ram[9159]  = 1;
  ram[9160]  = 1;
  ram[9161]  = 1;
  ram[9162]  = 1;
  ram[9163]  = 0;
  ram[9164]  = 1;
  ram[9165]  = 1;
  ram[9166]  = 1;
  ram[9167]  = 0;
  ram[9168]  = 1;
  ram[9169]  = 1;
  ram[9170]  = 1;
  ram[9171]  = 0;
  ram[9172]  = 1;
  ram[9173]  = 1;
  ram[9174]  = 1;
  ram[9175]  = 0;
  ram[9176]  = 0;
  ram[9177]  = 0;
  ram[9178]  = 0;
  ram[9179]  = 0;
  ram[9180]  = 0;
  ram[9181]  = 0;
  ram[9182]  = 0;
  ram[9183]  = 1;
  ram[9184]  = 1;
  ram[9185]  = 0;
  ram[9186]  = 1;
  ram[9187]  = 1;
  ram[9188]  = 1;
  ram[9189]  = 1;
  ram[9190]  = 1;
  ram[9191]  = 1;
  ram[9192]  = 0;
  ram[9193]  = 1;
  ram[9194]  = 1;
  ram[9195]  = 1;
  ram[9196]  = 1;
  ram[9197]  = 1;
  ram[9198]  = 1;
  ram[9199]  = 1;
  ram[9200]  = 1;
  ram[9201]  = 1;
  ram[9202]  = 1;
  ram[9203]  = 1;
  ram[9204]  = 1;
  ram[9205]  = 1;
  ram[9206]  = 1;
  ram[9207]  = 1;
  ram[9208]  = 1;
  ram[9209]  = 1;
  ram[9210]  = 1;
  ram[9211]  = 1;
  ram[9212]  = 1;
  ram[9213]  = 1;
  ram[9214]  = 1;
  ram[9215]  = 1;
  ram[9216]  = 1;
  ram[9217]  = 1;
  ram[9218]  = 1;
  ram[9219]  = 1;
  ram[9220]  = 1;
  ram[9221]  = 1;
  ram[9222]  = 1;
  ram[9223]  = 1;
  ram[9224]  = 1;
  ram[9225]  = 1;
  ram[9226]  = 1;
  ram[9227]  = 1;
  ram[9228]  = 1;
  ram[9229]  = 1;
  ram[9230]  = 1;
  ram[9231]  = 1;
  ram[9232]  = 1;
  ram[9233]  = 1;
  ram[9234]  = 1;
  ram[9235]  = 1;
  ram[9236]  = 1;
  ram[9237]  = 1;
  ram[9238]  = 1;
  ram[9239]  = 1;
  ram[9240]  = 1;
  ram[9241]  = 1;
  ram[9242]  = 1;
  ram[9243]  = 1;
  ram[9244]  = 1;
  ram[9245]  = 1;
  ram[9246]  = 1;
  ram[9247]  = 1;
  ram[9248]  = 1;
  ram[9249]  = 1;
  ram[9250]  = 1;
  ram[9251]  = 1;
  ram[9252]  = 1;
  ram[9253]  = 1;
  ram[9254]  = 1;
  ram[9255]  = 1;
  ram[9256]  = 1;
  ram[9257]  = 1;
  ram[9258]  = 1;
  ram[9259]  = 1;
  ram[9260]  = 1;
  ram[9261]  = 1;
  ram[9262]  = 1;
  ram[9263]  = 1;
  ram[9264]  = 1;
  ram[9265]  = 1;
  ram[9266]  = 1;
  ram[9267]  = 1;
  ram[9268]  = 1;
  ram[9269]  = 1;
  ram[9270]  = 1;
  ram[9271]  = 1;
  ram[9272]  = 1;
  ram[9273]  = 1;
  ram[9274]  = 1;
  ram[9275]  = 1;
  ram[9276]  = 1;
  ram[9277]  = 1;
  ram[9278]  = 1;
  ram[9279]  = 1;
  ram[9280]  = 1;
  ram[9281]  = 1;
  ram[9282]  = 1;
  ram[9283]  = 1;
  ram[9284]  = 1;
  ram[9285]  = 1;
  ram[9286]  = 1;
  ram[9287]  = 1;
  ram[9288]  = 1;
  ram[9289]  = 1;
  ram[9290]  = 1;
  ram[9291]  = 1;
  ram[9292]  = 1;
  ram[9293]  = 1;
  ram[9294]  = 1;
  ram[9295]  = 1;
  ram[9296]  = 1;
  ram[9297]  = 1;
  ram[9298]  = 1;
  ram[9299]  = 1;
  ram[9300]  = 1;
  ram[9301]  = 1;
  ram[9302]  = 1;
  ram[9303]  = 1;
  ram[9304]  = 1;
  ram[9305]  = 1;
  ram[9306]  = 1;
  ram[9307]  = 1;
  ram[9308]  = 1;
  ram[9309]  = 1;
  ram[9310]  = 1;
  ram[9311]  = 1;
  ram[9312]  = 1;
  ram[9313]  = 1;
  ram[9314]  = 1;
  ram[9315]  = 1;
  ram[9316]  = 1;
  ram[9317]  = 1;
  ram[9318]  = 1;
  ram[9319]  = 1;
  ram[9320]  = 1;
  ram[9321]  = 1;
  ram[9322]  = 1;
  ram[9323]  = 1;
  ram[9324]  = 1;
  ram[9325]  = 1;
  ram[9326]  = 1;
  ram[9327]  = 1;
  ram[9328]  = 1;
  ram[9329]  = 1;
  ram[9330]  = 1;
  ram[9331]  = 1;
  ram[9332]  = 1;
  ram[9333]  = 1;
  ram[9334]  = 1;
  ram[9335]  = 1;
  ram[9336]  = 1;
  ram[9337]  = 1;
  ram[9338]  = 1;
  ram[9339]  = 1;
  ram[9340]  = 1;
  ram[9341]  = 1;
  ram[9342]  = 1;
  ram[9343]  = 1;
  ram[9344]  = 1;
  ram[9345]  = 1;
  ram[9346]  = 1;
  ram[9347]  = 1;
  ram[9348]  = 1;
  ram[9349]  = 1;
  ram[9350]  = 1;
  ram[9351]  = 1;
  ram[9352]  = 1;
  ram[9353]  = 1;
  ram[9354]  = 1;
  ram[9355]  = 1;
  ram[9356]  = 1;
  ram[9357]  = 1;
  ram[9358]  = 1;
  ram[9359]  = 1;
  ram[9360]  = 1;
  ram[9361]  = 1;
  ram[9362]  = 1;
  ram[9363]  = 1;
  ram[9364]  = 1;
  ram[9365]  = 1;
  ram[9366]  = 1;
  ram[9367]  = 1;
  ram[9368]  = 1;
  ram[9369]  = 1;
  ram[9370]  = 1;
  ram[9371]  = 1;
  ram[9372]  = 1;
  ram[9373]  = 1;
  ram[9374]  = 1;
  ram[9375]  = 1;
  ram[9376]  = 1;
  ram[9377]  = 1;
  ram[9378]  = 1;
  ram[9379]  = 1;
  ram[9380]  = 1;
  ram[9381]  = 1;
  ram[9382]  = 1;
  ram[9383]  = 1;
  ram[9384]  = 1;
  ram[9385]  = 1;
  ram[9386]  = 1;
  ram[9387]  = 1;
  ram[9388]  = 1;
  ram[9389]  = 1;
  ram[9390]  = 1;
  ram[9391]  = 1;
  ram[9392]  = 1;
  ram[9393]  = 1;
  ram[9394]  = 1;
  ram[9395]  = 1;
  ram[9396]  = 1;
  ram[9397]  = 1;
  ram[9398]  = 1;
  ram[9399]  = 1;
  ram[9400]  = 0;
  ram[9401]  = 1;
  ram[9402]  = 1;
  ram[9403]  = 1;
  ram[9404]  = 1;
  ram[9405]  = 1;
  ram[9406]  = 1;
  ram[9407]  = 1;
  ram[9408]  = 1;
  ram[9409]  = 0;
  ram[9410]  = 1;
  ram[9411]  = 1;
  ram[9412]  = 1;
  ram[9413]  = 0;
  ram[9414]  = 0;
  ram[9415]  = 1;
  ram[9416]  = 1;
  ram[9417]  = 1;
  ram[9418]  = 0;
  ram[9419]  = 1;
  ram[9420]  = 1;
  ram[9421]  = 1;
  ram[9422]  = 0;
  ram[9423]  = 0;
  ram[9424]  = 1;
  ram[9425]  = 1;
  ram[9426]  = 1;
  ram[9427]  = 1;
  ram[9428]  = 0;
  ram[9429]  = 1;
  ram[9430]  = 1;
  ram[9431]  = 1;
  ram[9432]  = 1;
  ram[9433]  = 1;
  ram[9434]  = 0;
  ram[9435]  = 1;
  ram[9436]  = 1;
  ram[9437]  = 0;
  ram[9438]  = 0;
  ram[9439]  = 1;
  ram[9440]  = 1;
  ram[9441]  = 1;
  ram[9442]  = 1;
  ram[9443]  = 1;
  ram[9444]  = 1;
  ram[9445]  = 1;
  ram[9446]  = 1;
  ram[9447]  = 1;
  ram[9448]  = 1;
  ram[9449]  = 1;
  ram[9450]  = 1;
  ram[9451]  = 1;
  ram[9452]  = 0;
  ram[9453]  = 0;
  ram[9454]  = 1;
  ram[9455]  = 1;
  ram[9456]  = 1;
  ram[9457]  = 1;
  ram[9458]  = 1;
  ram[9459]  = 1;
  ram[9460]  = 1;
  ram[9461]  = 1;
  ram[9462]  = 1;
  ram[9463]  = 0;
  ram[9464]  = 1;
  ram[9465]  = 1;
  ram[9466]  = 1;
  ram[9467]  = 0;
  ram[9468]  = 1;
  ram[9469]  = 1;
  ram[9470]  = 0;
  ram[9471]  = 0;
  ram[9472]  = 1;
  ram[9473]  = 1;
  ram[9474]  = 1;
  ram[9475]  = 0;
  ram[9476]  = 1;
  ram[9477]  = 1;
  ram[9478]  = 1;
  ram[9479]  = 1;
  ram[9480]  = 1;
  ram[9481]  = 1;
  ram[9482]  = 1;
  ram[9483]  = 1;
  ram[9484]  = 1;
  ram[9485]  = 0;
  ram[9486]  = 1;
  ram[9487]  = 1;
  ram[9488]  = 1;
  ram[9489]  = 1;
  ram[9490]  = 1;
  ram[9491]  = 1;
  ram[9492]  = 0;
  ram[9493]  = 1;
  ram[9494]  = 1;
  ram[9495]  = 1;
  ram[9496]  = 1;
  ram[9497]  = 1;
  ram[9498]  = 1;
  ram[9499]  = 1;
  ram[9500]  = 1;
  ram[9501]  = 1;
  ram[9502]  = 1;
  ram[9503]  = 1;
  ram[9504]  = 1;
  ram[9505]  = 1;
  ram[9506]  = 1;
  ram[9507]  = 1;
  ram[9508]  = 1;
  ram[9509]  = 1;
  ram[9510]  = 1;
  ram[9511]  = 1;
  ram[9512]  = 1;
  ram[9513]  = 1;
  ram[9514]  = 1;
  ram[9515]  = 1;
  ram[9516]  = 1;
  ram[9517]  = 1;
  ram[9518]  = 1;
  ram[9519]  = 1;
  ram[9520]  = 1;
  ram[9521]  = 1;
  ram[9522]  = 1;
  ram[9523]  = 1;
  ram[9524]  = 1;
  ram[9525]  = 1;
  ram[9526]  = 1;
  ram[9527]  = 1;
  ram[9528]  = 1;
  ram[9529]  = 1;
  ram[9530]  = 1;
  ram[9531]  = 1;
  ram[9532]  = 1;
  ram[9533]  = 1;
  ram[9534]  = 1;
  ram[9535]  = 1;
  ram[9536]  = 1;
  ram[9537]  = 1;
  ram[9538]  = 1;
  ram[9539]  = 1;
  ram[9540]  = 1;
  ram[9541]  = 1;
  ram[9542]  = 1;
  ram[9543]  = 1;
  ram[9544]  = 1;
  ram[9545]  = 1;
  ram[9546]  = 1;
  ram[9547]  = 1;
  ram[9548]  = 1;
  ram[9549]  = 1;
  ram[9550]  = 1;
  ram[9551]  = 1;
  ram[9552]  = 1;
  ram[9553]  = 1;
  ram[9554]  = 1;
  ram[9555]  = 1;
  ram[9556]  = 1;
  ram[9557]  = 1;
  ram[9558]  = 1;
  ram[9559]  = 1;
  ram[9560]  = 1;
  ram[9561]  = 1;
  ram[9562]  = 1;
  ram[9563]  = 1;
  ram[9564]  = 1;
  ram[9565]  = 1;
  ram[9566]  = 1;
  ram[9567]  = 1;
  ram[9568]  = 1;
  ram[9569]  = 1;
  ram[9570]  = 1;
  ram[9571]  = 1;
  ram[9572]  = 1;
  ram[9573]  = 1;
  ram[9574]  = 1;
  ram[9575]  = 1;
  ram[9576]  = 1;
  ram[9577]  = 1;
  ram[9578]  = 1;
  ram[9579]  = 1;
  ram[9580]  = 1;
  ram[9581]  = 1;
  ram[9582]  = 1;
  ram[9583]  = 1;
  ram[9584]  = 1;
  ram[9585]  = 1;
  ram[9586]  = 1;
  ram[9587]  = 1;
  ram[9588]  = 1;
  ram[9589]  = 1;
  ram[9590]  = 1;
  ram[9591]  = 1;
  ram[9592]  = 1;
  ram[9593]  = 1;
  ram[9594]  = 1;
  ram[9595]  = 1;
  ram[9596]  = 1;
  ram[9597]  = 1;
  ram[9598]  = 1;
  ram[9599]  = 1;
  ram[9600]  = 1;
  ram[9601]  = 1;
  ram[9602]  = 1;
  ram[9603]  = 1;
  ram[9604]  = 1;
  ram[9605]  = 1;
  ram[9606]  = 1;
  ram[9607]  = 1;
  ram[9608]  = 1;
  ram[9609]  = 1;
  ram[9610]  = 1;
  ram[9611]  = 1;
  ram[9612]  = 1;
  ram[9613]  = 1;
  ram[9614]  = 1;
  ram[9615]  = 1;
  ram[9616]  = 1;
  ram[9617]  = 1;
  ram[9618]  = 1;
  ram[9619]  = 1;
  ram[9620]  = 1;
  ram[9621]  = 1;
  ram[9622]  = 1;
  ram[9623]  = 1;
  ram[9624]  = 1;
  ram[9625]  = 1;
  ram[9626]  = 1;
  ram[9627]  = 1;
  ram[9628]  = 1;
  ram[9629]  = 1;
  ram[9630]  = 1;
  ram[9631]  = 1;
  ram[9632]  = 1;
  ram[9633]  = 1;
  ram[9634]  = 1;
  ram[9635]  = 1;
  ram[9636]  = 1;
  ram[9637]  = 1;
  ram[9638]  = 1;
  ram[9639]  = 1;
  ram[9640]  = 1;
  ram[9641]  = 1;
  ram[9642]  = 1;
  ram[9643]  = 1;
  ram[9644]  = 1;
  ram[9645]  = 1;
  ram[9646]  = 1;
  ram[9647]  = 1;
  ram[9648]  = 1;
  ram[9649]  = 1;
  ram[9650]  = 1;
  ram[9651]  = 1;
  ram[9652]  = 1;
  ram[9653]  = 1;
  ram[9654]  = 1;
  ram[9655]  = 1;
  ram[9656]  = 1;
  ram[9657]  = 1;
  ram[9658]  = 1;
  ram[9659]  = 1;
  ram[9660]  = 1;
  ram[9661]  = 1;
  ram[9662]  = 1;
  ram[9663]  = 1;
  ram[9664]  = 1;
  ram[9665]  = 1;
  ram[9666]  = 1;
  ram[9667]  = 1;
  ram[9668]  = 1;
  ram[9669]  = 1;
  ram[9670]  = 1;
  ram[9671]  = 1;
  ram[9672]  = 1;
  ram[9673]  = 1;
  ram[9674]  = 1;
  ram[9675]  = 1;
  ram[9676]  = 1;
  ram[9677]  = 1;
  ram[9678]  = 1;
  ram[9679]  = 1;
  ram[9680]  = 1;
  ram[9681]  = 1;
  ram[9682]  = 1;
  ram[9683]  = 1;
  ram[9684]  = 1;
  ram[9685]  = 1;
  ram[9686]  = 1;
  ram[9687]  = 1;
  ram[9688]  = 1;
  ram[9689]  = 1;
  ram[9690]  = 1;
  ram[9691]  = 1;
  ram[9692]  = 1;
  ram[9693]  = 1;
  ram[9694]  = 1;
  ram[9695]  = 1;
  ram[9696]  = 1;
  ram[9697]  = 1;
  ram[9698]  = 1;
  ram[9699]  = 1;
  ram[9700]  = 0;
  ram[9701]  = 0;
  ram[9702]  = 1;
  ram[9703]  = 1;
  ram[9704]  = 1;
  ram[9705]  = 1;
  ram[9706]  = 1;
  ram[9707]  = 1;
  ram[9708]  = 1;
  ram[9709]  = 0;
  ram[9710]  = 1;
  ram[9711]  = 1;
  ram[9712]  = 1;
  ram[9713]  = 0;
  ram[9714]  = 1;
  ram[9715]  = 1;
  ram[9716]  = 1;
  ram[9717]  = 1;
  ram[9718]  = 0;
  ram[9719]  = 1;
  ram[9720]  = 1;
  ram[9721]  = 1;
  ram[9722]  = 0;
  ram[9723]  = 0;
  ram[9724]  = 1;
  ram[9725]  = 1;
  ram[9726]  = 1;
  ram[9727]  = 1;
  ram[9728]  = 0;
  ram[9729]  = 1;
  ram[9730]  = 1;
  ram[9731]  = 1;
  ram[9732]  = 1;
  ram[9733]  = 1;
  ram[9734]  = 0;
  ram[9735]  = 1;
  ram[9736]  = 1;
  ram[9737]  = 0;
  ram[9738]  = 0;
  ram[9739]  = 1;
  ram[9740]  = 1;
  ram[9741]  = 1;
  ram[9742]  = 1;
  ram[9743]  = 1;
  ram[9744]  = 1;
  ram[9745]  = 1;
  ram[9746]  = 1;
  ram[9747]  = 1;
  ram[9748]  = 1;
  ram[9749]  = 1;
  ram[9750]  = 1;
  ram[9751]  = 1;
  ram[9752]  = 0;
  ram[9753]  = 0;
  ram[9754]  = 1;
  ram[9755]  = 1;
  ram[9756]  = 1;
  ram[9757]  = 1;
  ram[9758]  = 1;
  ram[9759]  = 1;
  ram[9760]  = 1;
  ram[9761]  = 1;
  ram[9762]  = 0;
  ram[9763]  = 0;
  ram[9764]  = 1;
  ram[9765]  = 1;
  ram[9766]  = 1;
  ram[9767]  = 0;
  ram[9768]  = 1;
  ram[9769]  = 1;
  ram[9770]  = 0;
  ram[9771]  = 1;
  ram[9772]  = 1;
  ram[9773]  = 1;
  ram[9774]  = 1;
  ram[9775]  = 0;
  ram[9776]  = 1;
  ram[9777]  = 1;
  ram[9778]  = 1;
  ram[9779]  = 1;
  ram[9780]  = 1;
  ram[9781]  = 1;
  ram[9782]  = 1;
  ram[9783]  = 1;
  ram[9784]  = 1;
  ram[9785]  = 0;
  ram[9786]  = 1;
  ram[9787]  = 1;
  ram[9788]  = 1;
  ram[9789]  = 1;
  ram[9790]  = 1;
  ram[9791]  = 1;
  ram[9792]  = 0;
  ram[9793]  = 1;
  ram[9794]  = 1;
  ram[9795]  = 1;
  ram[9796]  = 1;
  ram[9797]  = 1;
  ram[9798]  = 1;
  ram[9799]  = 1;
  ram[9800]  = 1;
  ram[9801]  = 1;
  ram[9802]  = 1;
  ram[9803]  = 1;
  ram[9804]  = 1;
  ram[9805]  = 1;
  ram[9806]  = 1;
  ram[9807]  = 1;
  ram[9808]  = 1;
  ram[9809]  = 1;
  ram[9810]  = 1;
  ram[9811]  = 1;
  ram[9812]  = 1;
  ram[9813]  = 1;
  ram[9814]  = 1;
  ram[9815]  = 1;
  ram[9816]  = 1;
  ram[9817]  = 1;
  ram[9818]  = 1;
  ram[9819]  = 1;
  ram[9820]  = 1;
  ram[9821]  = 1;
  ram[9822]  = 1;
  ram[9823]  = 1;
  ram[9824]  = 1;
  ram[9825]  = 1;
  ram[9826]  = 1;
  ram[9827]  = 1;
  ram[9828]  = 1;
  ram[9829]  = 1;
  ram[9830]  = 1;
  ram[9831]  = 1;
  ram[9832]  = 1;
  ram[9833]  = 1;
  ram[9834]  = 1;
  ram[9835]  = 1;
  ram[9836]  = 1;
  ram[9837]  = 1;
  ram[9838]  = 1;
  ram[9839]  = 1;
  ram[9840]  = 1;
  ram[9841]  = 1;
  ram[9842]  = 1;
  ram[9843]  = 1;
  ram[9844]  = 1;
  ram[9845]  = 1;
  ram[9846]  = 1;
  ram[9847]  = 1;
  ram[9848]  = 1;
  ram[9849]  = 1;
  ram[9850]  = 1;
  ram[9851]  = 1;
  ram[9852]  = 1;
  ram[9853]  = 1;
  ram[9854]  = 1;
  ram[9855]  = 1;
  ram[9856]  = 1;
  ram[9857]  = 1;
  ram[9858]  = 1;
  ram[9859]  = 1;
  ram[9860]  = 1;
  ram[9861]  = 1;
  ram[9862]  = 1;
  ram[9863]  = 1;
  ram[9864]  = 1;
  ram[9865]  = 1;
  ram[9866]  = 1;
  ram[9867]  = 1;
  ram[9868]  = 1;
  ram[9869]  = 1;
  ram[9870]  = 1;
  ram[9871]  = 1;
  ram[9872]  = 1;
  ram[9873]  = 1;
  ram[9874]  = 1;
  ram[9875]  = 1;
  ram[9876]  = 1;
  ram[9877]  = 1;
  ram[9878]  = 1;
  ram[9879]  = 1;
  ram[9880]  = 1;
  ram[9881]  = 1;
  ram[9882]  = 1;
  ram[9883]  = 1;
  ram[9884]  = 1;
  ram[9885]  = 1;
  ram[9886]  = 1;
  ram[9887]  = 1;
  ram[9888]  = 1;
  ram[9889]  = 1;
  ram[9890]  = 1;
  ram[9891]  = 1;
  ram[9892]  = 1;
  ram[9893]  = 1;
  ram[9894]  = 1;
  ram[9895]  = 1;
  ram[9896]  = 1;
  ram[9897]  = 1;
  ram[9898]  = 1;
  ram[9899]  = 1;
  ram[9900]  = 1;
  ram[9901]  = 1;
  ram[9902]  = 1;
  ram[9903]  = 1;
  ram[9904]  = 1;
  ram[9905]  = 1;
  ram[9906]  = 1;
  ram[9907]  = 1;
  ram[9908]  = 1;
  ram[9909]  = 1;
  ram[9910]  = 1;
  ram[9911]  = 1;
  ram[9912]  = 1;
  ram[9913]  = 1;
  ram[9914]  = 1;
  ram[9915]  = 1;
  ram[9916]  = 1;
  ram[9917]  = 1;
  ram[9918]  = 1;
  ram[9919]  = 1;
  ram[9920]  = 1;
  ram[9921]  = 1;
  ram[9922]  = 1;
  ram[9923]  = 1;
  ram[9924]  = 1;
  ram[9925]  = 1;
  ram[9926]  = 1;
  ram[9927]  = 1;
  ram[9928]  = 1;
  ram[9929]  = 1;
  ram[9930]  = 1;
  ram[9931]  = 1;
  ram[9932]  = 1;
  ram[9933]  = 1;
  ram[9934]  = 1;
  ram[9935]  = 1;
  ram[9936]  = 1;
  ram[9937]  = 1;
  ram[9938]  = 1;
  ram[9939]  = 1;
  ram[9940]  = 1;
  ram[9941]  = 1;
  ram[9942]  = 1;
  ram[9943]  = 1;
  ram[9944]  = 1;
  ram[9945]  = 1;
  ram[9946]  = 1;
  ram[9947]  = 1;
  ram[9948]  = 1;
  ram[9949]  = 1;
  ram[9950]  = 1;
  ram[9951]  = 1;
  ram[9952]  = 1;
  ram[9953]  = 1;
  ram[9954]  = 1;
  ram[9955]  = 1;
  ram[9956]  = 1;
  ram[9957]  = 1;
  ram[9958]  = 1;
  ram[9959]  = 1;
  ram[9960]  = 1;
  ram[9961]  = 1;
  ram[9962]  = 1;
  ram[9963]  = 1;
  ram[9964]  = 1;
  ram[9965]  = 1;
  ram[9966]  = 1;
  ram[9967]  = 1;
  ram[9968]  = 1;
  ram[9969]  = 1;
  ram[9970]  = 1;
  ram[9971]  = 1;
  ram[9972]  = 1;
  ram[9973]  = 1;
  ram[9974]  = 1;
  ram[9975]  = 1;
  ram[9976]  = 1;
  ram[9977]  = 1;
  ram[9978]  = 1;
  ram[9979]  = 1;
  ram[9980]  = 1;
  ram[9981]  = 1;
  ram[9982]  = 1;
  ram[9983]  = 1;
  ram[9984]  = 1;
  ram[9985]  = 1;
  ram[9986]  = 1;
  ram[9987]  = 1;
  ram[9988]  = 1;
  ram[9989]  = 1;
  ram[9990]  = 1;
  ram[9991]  = 1;
  ram[9992]  = 1;
  ram[9993]  = 1;
  ram[9994]  = 1;
  ram[9995]  = 1;
  ram[9996]  = 1;
  ram[9997]  = 1;
  ram[9998]  = 1;
  ram[9999]  = 1;
  ram[10000]  = 0;
  ram[10001]  = 0;
  ram[10002]  = 1;
  ram[10003]  = 1;
  ram[10004]  = 1;
  ram[10005]  = 1;
  ram[10006]  = 1;
  ram[10007]  = 1;
  ram[10008]  = 1;
  ram[10009]  = 0;
  ram[10010]  = 1;
  ram[10011]  = 1;
  ram[10012]  = 0;
  ram[10013]  = 0;
  ram[10014]  = 1;
  ram[10015]  = 1;
  ram[10016]  = 1;
  ram[10017]  = 1;
  ram[10018]  = 0;
  ram[10019]  = 1;
  ram[10020]  = 1;
  ram[10021]  = 1;
  ram[10022]  = 0;
  ram[10023]  = 0;
  ram[10024]  = 1;
  ram[10025]  = 1;
  ram[10026]  = 1;
  ram[10027]  = 1;
  ram[10028]  = 0;
  ram[10029]  = 1;
  ram[10030]  = 1;
  ram[10031]  = 1;
  ram[10032]  = 1;
  ram[10033]  = 1;
  ram[10034]  = 0;
  ram[10035]  = 1;
  ram[10036]  = 1;
  ram[10037]  = 0;
  ram[10038]  = 0;
  ram[10039]  = 1;
  ram[10040]  = 1;
  ram[10041]  = 1;
  ram[10042]  = 1;
  ram[10043]  = 1;
  ram[10044]  = 1;
  ram[10045]  = 1;
  ram[10046]  = 1;
  ram[10047]  = 1;
  ram[10048]  = 1;
  ram[10049]  = 1;
  ram[10050]  = 1;
  ram[10051]  = 1;
  ram[10052]  = 1;
  ram[10053]  = 0;
  ram[10054]  = 1;
  ram[10055]  = 1;
  ram[10056]  = 1;
  ram[10057]  = 1;
  ram[10058]  = 1;
  ram[10059]  = 1;
  ram[10060]  = 1;
  ram[10061]  = 1;
  ram[10062]  = 0;
  ram[10063]  = 0;
  ram[10064]  = 1;
  ram[10065]  = 1;
  ram[10066]  = 1;
  ram[10067]  = 0;
  ram[10068]  = 0;
  ram[10069]  = 1;
  ram[10070]  = 0;
  ram[10071]  = 1;
  ram[10072]  = 1;
  ram[10073]  = 1;
  ram[10074]  = 1;
  ram[10075]  = 0;
  ram[10076]  = 1;
  ram[10077]  = 1;
  ram[10078]  = 1;
  ram[10079]  = 1;
  ram[10080]  = 1;
  ram[10081]  = 1;
  ram[10082]  = 1;
  ram[10083]  = 1;
  ram[10084]  = 1;
  ram[10085]  = 0;
  ram[10086]  = 1;
  ram[10087]  = 1;
  ram[10088]  = 1;
  ram[10089]  = 1;
  ram[10090]  = 1;
  ram[10091]  = 1;
  ram[10092]  = 1;
  ram[10093]  = 1;
  ram[10094]  = 1;
  ram[10095]  = 1;
  ram[10096]  = 1;
  ram[10097]  = 1;
  ram[10098]  = 1;
  ram[10099]  = 1;
  ram[10100]  = 1;
  ram[10101]  = 1;
  ram[10102]  = 1;
  ram[10103]  = 1;
  ram[10104]  = 1;
  ram[10105]  = 1;
  ram[10106]  = 1;
  ram[10107]  = 1;
  ram[10108]  = 1;
  ram[10109]  = 1;
  ram[10110]  = 1;
  ram[10111]  = 1;
  ram[10112]  = 1;
  ram[10113]  = 1;
  ram[10114]  = 1;
  ram[10115]  = 1;
  ram[10116]  = 1;
  ram[10117]  = 1;
  ram[10118]  = 1;
  ram[10119]  = 1;
  ram[10120]  = 1;
  ram[10121]  = 1;
  ram[10122]  = 1;
  ram[10123]  = 1;
  ram[10124]  = 1;
  ram[10125]  = 1;
  ram[10126]  = 1;
  ram[10127]  = 1;
  ram[10128]  = 1;
  ram[10129]  = 1;
  ram[10130]  = 1;
  ram[10131]  = 1;
  ram[10132]  = 1;
  ram[10133]  = 1;
  ram[10134]  = 1;
  ram[10135]  = 1;
  ram[10136]  = 1;
  ram[10137]  = 1;
  ram[10138]  = 1;
  ram[10139]  = 1;
  ram[10140]  = 1;
  ram[10141]  = 1;
  ram[10142]  = 1;
  ram[10143]  = 1;
  ram[10144]  = 1;
  ram[10145]  = 1;
  ram[10146]  = 1;
  ram[10147]  = 1;
  ram[10148]  = 1;
  ram[10149]  = 1;
  ram[10150]  = 1;
  ram[10151]  = 1;
  ram[10152]  = 1;
  ram[10153]  = 1;
  ram[10154]  = 1;
  ram[10155]  = 1;
  ram[10156]  = 1;
  ram[10157]  = 1;
  ram[10158]  = 1;
  ram[10159]  = 1;
  ram[10160]  = 1;
  ram[10161]  = 1;
  ram[10162]  = 1;
  ram[10163]  = 1;
  ram[10164]  = 1;
  ram[10165]  = 1;
  ram[10166]  = 1;
  ram[10167]  = 1;
  ram[10168]  = 1;
  ram[10169]  = 1;
  ram[10170]  = 1;
  ram[10171]  = 1;
  ram[10172]  = 1;
  ram[10173]  = 1;
  ram[10174]  = 1;
  ram[10175]  = 1;
  ram[10176]  = 1;
  ram[10177]  = 1;
  ram[10178]  = 1;
  ram[10179]  = 1;
  ram[10180]  = 1;
  ram[10181]  = 1;
  ram[10182]  = 1;
  ram[10183]  = 1;
  ram[10184]  = 1;
  ram[10185]  = 1;
  ram[10186]  = 1;
  ram[10187]  = 1;
  ram[10188]  = 1;
  ram[10189]  = 1;
  ram[10190]  = 1;
  ram[10191]  = 1;
  ram[10192]  = 1;
  ram[10193]  = 1;
  ram[10194]  = 1;
  ram[10195]  = 1;
  ram[10196]  = 1;
  ram[10197]  = 1;
  ram[10198]  = 1;
  ram[10199]  = 1;
  ram[10200]  = 1;
  ram[10201]  = 1;
  ram[10202]  = 1;
  ram[10203]  = 1;
  ram[10204]  = 1;
  ram[10205]  = 1;
  ram[10206]  = 1;
  ram[10207]  = 1;
  ram[10208]  = 1;
  ram[10209]  = 1;
  ram[10210]  = 1;
  ram[10211]  = 1;
  ram[10212]  = 1;
  ram[10213]  = 1;
  ram[10214]  = 1;
  ram[10215]  = 1;
  ram[10216]  = 1;
  ram[10217]  = 1;
  ram[10218]  = 1;
  ram[10219]  = 1;
  ram[10220]  = 1;
  ram[10221]  = 1;
  ram[10222]  = 1;
  ram[10223]  = 1;
  ram[10224]  = 1;
  ram[10225]  = 1;
  ram[10226]  = 1;
  ram[10227]  = 1;
  ram[10228]  = 1;
  ram[10229]  = 1;
  ram[10230]  = 1;
  ram[10231]  = 1;
  ram[10232]  = 1;
  ram[10233]  = 1;
  ram[10234]  = 1;
  ram[10235]  = 1;
  ram[10236]  = 1;
  ram[10237]  = 1;
  ram[10238]  = 1;
  ram[10239]  = 1;
  ram[10240]  = 1;
  ram[10241]  = 1;
  ram[10242]  = 1;
  ram[10243]  = 1;
  ram[10244]  = 1;
  ram[10245]  = 1;
  ram[10246]  = 1;
  ram[10247]  = 1;
  ram[10248]  = 1;
  ram[10249]  = 1;
  ram[10250]  = 1;
  ram[10251]  = 1;
  ram[10252]  = 1;
  ram[10253]  = 1;
  ram[10254]  = 1;
  ram[10255]  = 1;
  ram[10256]  = 1;
  ram[10257]  = 1;
  ram[10258]  = 1;
  ram[10259]  = 1;
  ram[10260]  = 1;
  ram[10261]  = 1;
  ram[10262]  = 1;
  ram[10263]  = 1;
  ram[10264]  = 1;
  ram[10265]  = 1;
  ram[10266]  = 1;
  ram[10267]  = 1;
  ram[10268]  = 1;
  ram[10269]  = 1;
  ram[10270]  = 1;
  ram[10271]  = 1;
  ram[10272]  = 1;
  ram[10273]  = 1;
  ram[10274]  = 1;
  ram[10275]  = 1;
  ram[10276]  = 1;
  ram[10277]  = 1;
  ram[10278]  = 1;
  ram[10279]  = 1;
  ram[10280]  = 1;
  ram[10281]  = 1;
  ram[10282]  = 1;
  ram[10283]  = 1;
  ram[10284]  = 1;
  ram[10285]  = 1;
  ram[10286]  = 1;
  ram[10287]  = 1;
  ram[10288]  = 1;
  ram[10289]  = 1;
  ram[10290]  = 1;
  ram[10291]  = 1;
  ram[10292]  = 1;
  ram[10293]  = 1;
  ram[10294]  = 1;
  ram[10295]  = 1;
  ram[10296]  = 1;
  ram[10297]  = 1;
  ram[10298]  = 1;
  ram[10299]  = 1;
  ram[10300]  = 1;
  ram[10301]  = 0;
  ram[10302]  = 1;
  ram[10303]  = 1;
  ram[10304]  = 1;
  ram[10305]  = 1;
  ram[10306]  = 1;
  ram[10307]  = 1;
  ram[10308]  = 1;
  ram[10309]  = 0;
  ram[10310]  = 1;
  ram[10311]  = 1;
  ram[10312]  = 0;
  ram[10313]  = 0;
  ram[10314]  = 1;
  ram[10315]  = 1;
  ram[10316]  = 1;
  ram[10317]  = 1;
  ram[10318]  = 0;
  ram[10319]  = 1;
  ram[10320]  = 1;
  ram[10321]  = 1;
  ram[10322]  = 0;
  ram[10323]  = 0;
  ram[10324]  = 1;
  ram[10325]  = 1;
  ram[10326]  = 1;
  ram[10327]  = 1;
  ram[10328]  = 0;
  ram[10329]  = 1;
  ram[10330]  = 1;
  ram[10331]  = 1;
  ram[10332]  = 1;
  ram[10333]  = 1;
  ram[10334]  = 0;
  ram[10335]  = 1;
  ram[10336]  = 1;
  ram[10337]  = 1;
  ram[10338]  = 0;
  ram[10339]  = 1;
  ram[10340]  = 1;
  ram[10341]  = 1;
  ram[10342]  = 1;
  ram[10343]  = 1;
  ram[10344]  = 1;
  ram[10345]  = 1;
  ram[10346]  = 1;
  ram[10347]  = 1;
  ram[10348]  = 1;
  ram[10349]  = 1;
  ram[10350]  = 1;
  ram[10351]  = 1;
  ram[10352]  = 1;
  ram[10353]  = 0;
  ram[10354]  = 1;
  ram[10355]  = 1;
  ram[10356]  = 1;
  ram[10357]  = 1;
  ram[10358]  = 1;
  ram[10359]  = 1;
  ram[10360]  = 1;
  ram[10361]  = 1;
  ram[10362]  = 0;
  ram[10363]  = 1;
  ram[10364]  = 1;
  ram[10365]  = 1;
  ram[10366]  = 1;
  ram[10367]  = 1;
  ram[10368]  = 0;
  ram[10369]  = 1;
  ram[10370]  = 0;
  ram[10371]  = 1;
  ram[10372]  = 1;
  ram[10373]  = 1;
  ram[10374]  = 1;
  ram[10375]  = 0;
  ram[10376]  = 1;
  ram[10377]  = 1;
  ram[10378]  = 1;
  ram[10379]  = 1;
  ram[10380]  = 1;
  ram[10381]  = 1;
  ram[10382]  = 1;
  ram[10383]  = 1;
  ram[10384]  = 1;
  ram[10385]  = 0;
  ram[10386]  = 1;
  ram[10387]  = 1;
  ram[10388]  = 1;
  ram[10389]  = 1;
  ram[10390]  = 1;
  ram[10391]  = 1;
  ram[10392]  = 1;
  ram[10393]  = 1;
  ram[10394]  = 1;
  ram[10395]  = 1;
  ram[10396]  = 1;
  ram[10397]  = 1;
  ram[10398]  = 1;
  ram[10399]  = 1;
  ram[10400]  = 1;
  ram[10401]  = 1;
  ram[10402]  = 1;
  ram[10403]  = 1;
  ram[10404]  = 1;
  ram[10405]  = 1;
  ram[10406]  = 1;
  ram[10407]  = 1;
  ram[10408]  = 1;
  ram[10409]  = 1;
  ram[10410]  = 1;
  ram[10411]  = 1;
  ram[10412]  = 1;
  ram[10413]  = 1;
  ram[10414]  = 1;
  ram[10415]  = 1;
  ram[10416]  = 1;
  ram[10417]  = 1;
  ram[10418]  = 1;
  ram[10419]  = 1;
  ram[10420]  = 1;
  ram[10421]  = 1;
  ram[10422]  = 1;
  ram[10423]  = 1;
  ram[10424]  = 1;
  ram[10425]  = 1;
  ram[10426]  = 1;
  ram[10427]  = 1;
  ram[10428]  = 1;
  ram[10429]  = 1;
  ram[10430]  = 1;
  ram[10431]  = 1;
  ram[10432]  = 1;
  ram[10433]  = 1;
  ram[10434]  = 1;
  ram[10435]  = 1;
  ram[10436]  = 1;
  ram[10437]  = 1;
  ram[10438]  = 1;
  ram[10439]  = 1;
  ram[10440]  = 1;
  ram[10441]  = 1;
  ram[10442]  = 1;
  ram[10443]  = 1;
  ram[10444]  = 1;
  ram[10445]  = 1;
  ram[10446]  = 1;
  ram[10447]  = 1;
  ram[10448]  = 1;
  ram[10449]  = 1;
  ram[10450]  = 1;
  ram[10451]  = 1;
  ram[10452]  = 1;
  ram[10453]  = 1;
  ram[10454]  = 1;
  ram[10455]  = 1;
  ram[10456]  = 1;
  ram[10457]  = 1;
  ram[10458]  = 1;
  ram[10459]  = 1;
  ram[10460]  = 1;
  ram[10461]  = 1;
  ram[10462]  = 1;
  ram[10463]  = 1;
  ram[10464]  = 1;
  ram[10465]  = 1;
  ram[10466]  = 1;
  ram[10467]  = 1;
  ram[10468]  = 1;
  ram[10469]  = 1;
  ram[10470]  = 1;
  ram[10471]  = 1;
  ram[10472]  = 1;
  ram[10473]  = 1;
  ram[10474]  = 1;
  ram[10475]  = 1;
  ram[10476]  = 1;
  ram[10477]  = 1;
  ram[10478]  = 1;
  ram[10479]  = 1;
  ram[10480]  = 1;
  ram[10481]  = 1;
  ram[10482]  = 1;
  ram[10483]  = 1;
  ram[10484]  = 1;
  ram[10485]  = 1;
  ram[10486]  = 1;
  ram[10487]  = 1;
  ram[10488]  = 1;
  ram[10489]  = 1;
  ram[10490]  = 1;
  ram[10491]  = 1;
  ram[10492]  = 1;
  ram[10493]  = 1;
  ram[10494]  = 1;
  ram[10495]  = 1;
  ram[10496]  = 1;
  ram[10497]  = 1;
  ram[10498]  = 1;
  ram[10499]  = 1;
  ram[10500]  = 1;
  ram[10501]  = 1;
  ram[10502]  = 1;
  ram[10503]  = 1;
  ram[10504]  = 1;
  ram[10505]  = 1;
  ram[10506]  = 1;
  ram[10507]  = 1;
  ram[10508]  = 1;
  ram[10509]  = 1;
  ram[10510]  = 1;
  ram[10511]  = 1;
  ram[10512]  = 1;
  ram[10513]  = 1;
  ram[10514]  = 1;
  ram[10515]  = 1;
  ram[10516]  = 1;
  ram[10517]  = 1;
  ram[10518]  = 1;
  ram[10519]  = 1;
  ram[10520]  = 1;
  ram[10521]  = 1;
  ram[10522]  = 1;
  ram[10523]  = 1;
  ram[10524]  = 1;
  ram[10525]  = 1;
  ram[10526]  = 1;
  ram[10527]  = 1;
  ram[10528]  = 1;
  ram[10529]  = 1;
  ram[10530]  = 1;
  ram[10531]  = 1;
  ram[10532]  = 1;
  ram[10533]  = 1;
  ram[10534]  = 1;
  ram[10535]  = 1;
  ram[10536]  = 1;
  ram[10537]  = 1;
  ram[10538]  = 1;
  ram[10539]  = 1;
  ram[10540]  = 1;
  ram[10541]  = 1;
  ram[10542]  = 1;
  ram[10543]  = 1;
  ram[10544]  = 1;
  ram[10545]  = 1;
  ram[10546]  = 1;
  ram[10547]  = 1;
  ram[10548]  = 1;
  ram[10549]  = 1;
  ram[10550]  = 1;
  ram[10551]  = 1;
  ram[10552]  = 1;
  ram[10553]  = 1;
  ram[10554]  = 1;
  ram[10555]  = 1;
  ram[10556]  = 1;
  ram[10557]  = 1;
  ram[10558]  = 1;
  ram[10559]  = 1;
  ram[10560]  = 1;
  ram[10561]  = 1;
  ram[10562]  = 1;
  ram[10563]  = 1;
  ram[10564]  = 1;
  ram[10565]  = 1;
  ram[10566]  = 1;
  ram[10567]  = 1;
  ram[10568]  = 1;
  ram[10569]  = 1;
  ram[10570]  = 1;
  ram[10571]  = 1;
  ram[10572]  = 1;
  ram[10573]  = 1;
  ram[10574]  = 1;
  ram[10575]  = 1;
  ram[10576]  = 1;
  ram[10577]  = 1;
  ram[10578]  = 1;
  ram[10579]  = 1;
  ram[10580]  = 1;
  ram[10581]  = 1;
  ram[10582]  = 1;
  ram[10583]  = 1;
  ram[10584]  = 1;
  ram[10585]  = 1;
  ram[10586]  = 1;
  ram[10587]  = 1;
  ram[10588]  = 1;
  ram[10589]  = 1;
  ram[10590]  = 1;
  ram[10591]  = 1;
  ram[10592]  = 1;
  ram[10593]  = 1;
  ram[10594]  = 1;
  ram[10595]  = 1;
  ram[10596]  = 1;
  ram[10597]  = 1;
  ram[10598]  = 1;
  ram[10599]  = 1;
  ram[10600]  = 1;
  ram[10601]  = 0;
  ram[10602]  = 0;
  ram[10603]  = 1;
  ram[10604]  = 1;
  ram[10605]  = 1;
  ram[10606]  = 1;
  ram[10607]  = 1;
  ram[10608]  = 1;
  ram[10609]  = 0;
  ram[10610]  = 1;
  ram[10611]  = 1;
  ram[10612]  = 0;
  ram[10613]  = 0;
  ram[10614]  = 1;
  ram[10615]  = 1;
  ram[10616]  = 1;
  ram[10617]  = 1;
  ram[10618]  = 0;
  ram[10619]  = 1;
  ram[10620]  = 1;
  ram[10621]  = 1;
  ram[10622]  = 0;
  ram[10623]  = 0;
  ram[10624]  = 1;
  ram[10625]  = 1;
  ram[10626]  = 1;
  ram[10627]  = 1;
  ram[10628]  = 0;
  ram[10629]  = 1;
  ram[10630]  = 1;
  ram[10631]  = 1;
  ram[10632]  = 1;
  ram[10633]  = 1;
  ram[10634]  = 0;
  ram[10635]  = 1;
  ram[10636]  = 1;
  ram[10637]  = 1;
  ram[10638]  = 0;
  ram[10639]  = 1;
  ram[10640]  = 1;
  ram[10641]  = 1;
  ram[10642]  = 1;
  ram[10643]  = 1;
  ram[10644]  = 0;
  ram[10645]  = 1;
  ram[10646]  = 1;
  ram[10647]  = 1;
  ram[10648]  = 1;
  ram[10649]  = 1;
  ram[10650]  = 1;
  ram[10651]  = 1;
  ram[10652]  = 1;
  ram[10653]  = 0;
  ram[10654]  = 0;
  ram[10655]  = 1;
  ram[10656]  = 1;
  ram[10657]  = 1;
  ram[10658]  = 1;
  ram[10659]  = 1;
  ram[10660]  = 1;
  ram[10661]  = 0;
  ram[10662]  = 0;
  ram[10663]  = 1;
  ram[10664]  = 1;
  ram[10665]  = 1;
  ram[10666]  = 1;
  ram[10667]  = 1;
  ram[10668]  = 0;
  ram[10669]  = 1;
  ram[10670]  = 0;
  ram[10671]  = 1;
  ram[10672]  = 1;
  ram[10673]  = 1;
  ram[10674]  = 1;
  ram[10675]  = 0;
  ram[10676]  = 1;
  ram[10677]  = 1;
  ram[10678]  = 1;
  ram[10679]  = 1;
  ram[10680]  = 1;
  ram[10681]  = 0;
  ram[10682]  = 1;
  ram[10683]  = 1;
  ram[10684]  = 1;
  ram[10685]  = 0;
  ram[10686]  = 1;
  ram[10687]  = 1;
  ram[10688]  = 1;
  ram[10689]  = 1;
  ram[10690]  = 1;
  ram[10691]  = 1;
  ram[10692]  = 1;
  ram[10693]  = 1;
  ram[10694]  = 1;
  ram[10695]  = 1;
  ram[10696]  = 1;
  ram[10697]  = 1;
  ram[10698]  = 1;
  ram[10699]  = 1;
  ram[10700]  = 1;
  ram[10701]  = 1;
  ram[10702]  = 1;
  ram[10703]  = 1;
  ram[10704]  = 1;
  ram[10705]  = 1;
  ram[10706]  = 1;
  ram[10707]  = 1;
  ram[10708]  = 1;
  ram[10709]  = 1;
  ram[10710]  = 1;
  ram[10711]  = 1;
  ram[10712]  = 1;
  ram[10713]  = 1;
  ram[10714]  = 1;
  ram[10715]  = 1;
  ram[10716]  = 1;
  ram[10717]  = 1;
  ram[10718]  = 1;
  ram[10719]  = 1;
  ram[10720]  = 1;
  ram[10721]  = 1;
  ram[10722]  = 1;
  ram[10723]  = 1;
  ram[10724]  = 1;
  ram[10725]  = 1;
  ram[10726]  = 1;
  ram[10727]  = 1;
  ram[10728]  = 1;
  ram[10729]  = 1;
  ram[10730]  = 1;
  ram[10731]  = 1;
  ram[10732]  = 1;
  ram[10733]  = 1;
  ram[10734]  = 1;
  ram[10735]  = 1;
  ram[10736]  = 1;
  ram[10737]  = 1;
  ram[10738]  = 1;
  ram[10739]  = 1;
  ram[10740]  = 1;
  ram[10741]  = 1;
  ram[10742]  = 1;
  ram[10743]  = 1;
  ram[10744]  = 1;
  ram[10745]  = 1;
  ram[10746]  = 1;
  ram[10747]  = 1;
  ram[10748]  = 1;
  ram[10749]  = 1;
  ram[10750]  = 1;
  ram[10751]  = 1;
  ram[10752]  = 1;
  ram[10753]  = 1;
  ram[10754]  = 1;
  ram[10755]  = 1;
  ram[10756]  = 1;
  ram[10757]  = 1;
  ram[10758]  = 1;
  ram[10759]  = 1;
  ram[10760]  = 1;
  ram[10761]  = 1;
  ram[10762]  = 1;
  ram[10763]  = 1;
  ram[10764]  = 1;
  ram[10765]  = 1;
  ram[10766]  = 1;
  ram[10767]  = 1;
  ram[10768]  = 1;
  ram[10769]  = 1;
  ram[10770]  = 1;
  ram[10771]  = 1;
  ram[10772]  = 1;
  ram[10773]  = 1;
  ram[10774]  = 1;
  ram[10775]  = 1;
  ram[10776]  = 1;
  ram[10777]  = 1;
  ram[10778]  = 1;
  ram[10779]  = 1;
  ram[10780]  = 1;
  ram[10781]  = 1;
  ram[10782]  = 1;
  ram[10783]  = 1;
  ram[10784]  = 1;
  ram[10785]  = 1;
  ram[10786]  = 1;
  ram[10787]  = 1;
  ram[10788]  = 1;
  ram[10789]  = 1;
  ram[10790]  = 1;
  ram[10791]  = 1;
  ram[10792]  = 1;
  ram[10793]  = 1;
  ram[10794]  = 1;
  ram[10795]  = 1;
  ram[10796]  = 1;
  ram[10797]  = 1;
  ram[10798]  = 1;
  ram[10799]  = 1;
  ram[10800]  = 1;
  ram[10801]  = 1;
  ram[10802]  = 1;
  ram[10803]  = 1;
  ram[10804]  = 1;
  ram[10805]  = 1;
  ram[10806]  = 1;
  ram[10807]  = 1;
  ram[10808]  = 1;
  ram[10809]  = 1;
  ram[10810]  = 1;
  ram[10811]  = 1;
  ram[10812]  = 1;
  ram[10813]  = 1;
  ram[10814]  = 1;
  ram[10815]  = 1;
  ram[10816]  = 1;
  ram[10817]  = 1;
  ram[10818]  = 1;
  ram[10819]  = 1;
  ram[10820]  = 1;
  ram[10821]  = 1;
  ram[10822]  = 1;
  ram[10823]  = 1;
  ram[10824]  = 1;
  ram[10825]  = 1;
  ram[10826]  = 1;
  ram[10827]  = 1;
  ram[10828]  = 1;
  ram[10829]  = 1;
  ram[10830]  = 1;
  ram[10831]  = 1;
  ram[10832]  = 1;
  ram[10833]  = 1;
  ram[10834]  = 1;
  ram[10835]  = 1;
  ram[10836]  = 1;
  ram[10837]  = 1;
  ram[10838]  = 1;
  ram[10839]  = 1;
  ram[10840]  = 1;
  ram[10841]  = 1;
  ram[10842]  = 1;
  ram[10843]  = 1;
  ram[10844]  = 1;
  ram[10845]  = 1;
  ram[10846]  = 1;
  ram[10847]  = 1;
  ram[10848]  = 1;
  ram[10849]  = 1;
  ram[10850]  = 1;
  ram[10851]  = 1;
  ram[10852]  = 1;
  ram[10853]  = 1;
  ram[10854]  = 1;
  ram[10855]  = 1;
  ram[10856]  = 1;
  ram[10857]  = 1;
  ram[10858]  = 1;
  ram[10859]  = 1;
  ram[10860]  = 1;
  ram[10861]  = 1;
  ram[10862]  = 1;
  ram[10863]  = 1;
  ram[10864]  = 1;
  ram[10865]  = 1;
  ram[10866]  = 1;
  ram[10867]  = 1;
  ram[10868]  = 1;
  ram[10869]  = 1;
  ram[10870]  = 1;
  ram[10871]  = 1;
  ram[10872]  = 1;
  ram[10873]  = 1;
  ram[10874]  = 1;
  ram[10875]  = 1;
  ram[10876]  = 1;
  ram[10877]  = 1;
  ram[10878]  = 1;
  ram[10879]  = 1;
  ram[10880]  = 1;
  ram[10881]  = 1;
  ram[10882]  = 1;
  ram[10883]  = 1;
  ram[10884]  = 1;
  ram[10885]  = 1;
  ram[10886]  = 1;
  ram[10887]  = 1;
  ram[10888]  = 1;
  ram[10889]  = 1;
  ram[10890]  = 1;
  ram[10891]  = 1;
  ram[10892]  = 1;
  ram[10893]  = 1;
  ram[10894]  = 1;
  ram[10895]  = 1;
  ram[10896]  = 1;
  ram[10897]  = 1;
  ram[10898]  = 1;
  ram[10899]  = 1;
  ram[10900]  = 1;
  ram[10901]  = 1;
  ram[10902]  = 0;
  ram[10903]  = 1;
  ram[10904]  = 1;
  ram[10905]  = 1;
  ram[10906]  = 1;
  ram[10907]  = 1;
  ram[10908]  = 0;
  ram[10909]  = 0;
  ram[10910]  = 1;
  ram[10911]  = 1;
  ram[10912]  = 0;
  ram[10913]  = 0;
  ram[10914]  = 1;
  ram[10915]  = 1;
  ram[10916]  = 1;
  ram[10917]  = 0;
  ram[10918]  = 0;
  ram[10919]  = 1;
  ram[10920]  = 1;
  ram[10921]  = 1;
  ram[10922]  = 0;
  ram[10923]  = 0;
  ram[10924]  = 1;
  ram[10925]  = 1;
  ram[10926]  = 1;
  ram[10927]  = 1;
  ram[10928]  = 0;
  ram[10929]  = 1;
  ram[10930]  = 1;
  ram[10931]  = 1;
  ram[10932]  = 1;
  ram[10933]  = 1;
  ram[10934]  = 0;
  ram[10935]  = 1;
  ram[10936]  = 1;
  ram[10937]  = 1;
  ram[10938]  = 0;
  ram[10939]  = 0;
  ram[10940]  = 1;
  ram[10941]  = 1;
  ram[10942]  = 1;
  ram[10943]  = 0;
  ram[10944]  = 0;
  ram[10945]  = 1;
  ram[10946]  = 1;
  ram[10947]  = 1;
  ram[10948]  = 1;
  ram[10949]  = 1;
  ram[10950]  = 1;
  ram[10951]  = 1;
  ram[10952]  = 1;
  ram[10953]  = 1;
  ram[10954]  = 0;
  ram[10955]  = 1;
  ram[10956]  = 1;
  ram[10957]  = 1;
  ram[10958]  = 1;
  ram[10959]  = 1;
  ram[10960]  = 1;
  ram[10961]  = 0;
  ram[10962]  = 1;
  ram[10963]  = 1;
  ram[10964]  = 1;
  ram[10965]  = 1;
  ram[10966]  = 1;
  ram[10967]  = 1;
  ram[10968]  = 0;
  ram[10969]  = 0;
  ram[10970]  = 0;
  ram[10971]  = 1;
  ram[10972]  = 1;
  ram[10973]  = 1;
  ram[10974]  = 1;
  ram[10975]  = 0;
  ram[10976]  = 0;
  ram[10977]  = 1;
  ram[10978]  = 1;
  ram[10979]  = 1;
  ram[10980]  = 1;
  ram[10981]  = 0;
  ram[10982]  = 1;
  ram[10983]  = 1;
  ram[10984]  = 1;
  ram[10985]  = 0;
  ram[10986]  = 1;
  ram[10987]  = 1;
  ram[10988]  = 1;
  ram[10989]  = 1;
  ram[10990]  = 1;
  ram[10991]  = 1;
  ram[10992]  = 1;
  ram[10993]  = 1;
  ram[10994]  = 1;
  ram[10995]  = 1;
  ram[10996]  = 1;
  ram[10997]  = 1;
  ram[10998]  = 1;
  ram[10999]  = 1;
  ram[11000]  = 1;
  ram[11001]  = 1;
  ram[11002]  = 1;
  ram[11003]  = 1;
  ram[11004]  = 1;
  ram[11005]  = 1;
  ram[11006]  = 1;
  ram[11007]  = 1;
  ram[11008]  = 1;
  ram[11009]  = 1;
  ram[11010]  = 1;
  ram[11011]  = 1;
  ram[11012]  = 1;
  ram[11013]  = 1;
  ram[11014]  = 1;
  ram[11015]  = 1;
  ram[11016]  = 1;
  ram[11017]  = 1;
  ram[11018]  = 1;
  ram[11019]  = 1;
  ram[11020]  = 1;
  ram[11021]  = 1;
  ram[11022]  = 1;
  ram[11023]  = 1;
  ram[11024]  = 1;
  ram[11025]  = 1;
  ram[11026]  = 1;
  ram[11027]  = 1;
  ram[11028]  = 1;
  ram[11029]  = 1;
  ram[11030]  = 1;
  ram[11031]  = 1;
  ram[11032]  = 1;
  ram[11033]  = 1;
  ram[11034]  = 1;
  ram[11035]  = 1;
  ram[11036]  = 1;
  ram[11037]  = 1;
  ram[11038]  = 1;
  ram[11039]  = 1;
  ram[11040]  = 1;
  ram[11041]  = 1;
  ram[11042]  = 1;
  ram[11043]  = 1;
  ram[11044]  = 1;
  ram[11045]  = 1;
  ram[11046]  = 1;
  ram[11047]  = 1;
  ram[11048]  = 1;
  ram[11049]  = 1;
  ram[11050]  = 1;
  ram[11051]  = 1;
  ram[11052]  = 1;
  ram[11053]  = 1;
  ram[11054]  = 1;
  ram[11055]  = 1;
  ram[11056]  = 1;
  ram[11057]  = 1;
  ram[11058]  = 1;
  ram[11059]  = 1;
  ram[11060]  = 1;
  ram[11061]  = 1;
  ram[11062]  = 1;
  ram[11063]  = 1;
  ram[11064]  = 1;
  ram[11065]  = 1;
  ram[11066]  = 1;
  ram[11067]  = 1;
  ram[11068]  = 1;
  ram[11069]  = 1;
  ram[11070]  = 1;
  ram[11071]  = 1;
  ram[11072]  = 1;
  ram[11073]  = 1;
  ram[11074]  = 1;
  ram[11075]  = 1;
  ram[11076]  = 1;
  ram[11077]  = 1;
  ram[11078]  = 1;
  ram[11079]  = 1;
  ram[11080]  = 1;
  ram[11081]  = 1;
  ram[11082]  = 1;
  ram[11083]  = 1;
  ram[11084]  = 1;
  ram[11085]  = 1;
  ram[11086]  = 1;
  ram[11087]  = 1;
  ram[11088]  = 1;
  ram[11089]  = 1;
  ram[11090]  = 1;
  ram[11091]  = 1;
  ram[11092]  = 1;
  ram[11093]  = 1;
  ram[11094]  = 1;
  ram[11095]  = 1;
  ram[11096]  = 1;
  ram[11097]  = 1;
  ram[11098]  = 1;
  ram[11099]  = 1;
  ram[11100]  = 1;
  ram[11101]  = 1;
  ram[11102]  = 1;
  ram[11103]  = 1;
  ram[11104]  = 1;
  ram[11105]  = 1;
  ram[11106]  = 1;
  ram[11107]  = 1;
  ram[11108]  = 1;
  ram[11109]  = 1;
  ram[11110]  = 1;
  ram[11111]  = 1;
  ram[11112]  = 1;
  ram[11113]  = 1;
  ram[11114]  = 1;
  ram[11115]  = 1;
  ram[11116]  = 1;
  ram[11117]  = 1;
  ram[11118]  = 1;
  ram[11119]  = 1;
  ram[11120]  = 1;
  ram[11121]  = 1;
  ram[11122]  = 1;
  ram[11123]  = 1;
  ram[11124]  = 1;
  ram[11125]  = 1;
  ram[11126]  = 1;
  ram[11127]  = 1;
  ram[11128]  = 1;
  ram[11129]  = 1;
  ram[11130]  = 1;
  ram[11131]  = 1;
  ram[11132]  = 1;
  ram[11133]  = 1;
  ram[11134]  = 1;
  ram[11135]  = 1;
  ram[11136]  = 1;
  ram[11137]  = 1;
  ram[11138]  = 1;
  ram[11139]  = 1;
  ram[11140]  = 1;
  ram[11141]  = 1;
  ram[11142]  = 1;
  ram[11143]  = 1;
  ram[11144]  = 1;
  ram[11145]  = 1;
  ram[11146]  = 1;
  ram[11147]  = 1;
  ram[11148]  = 1;
  ram[11149]  = 1;
  ram[11150]  = 1;
  ram[11151]  = 1;
  ram[11152]  = 1;
  ram[11153]  = 1;
  ram[11154]  = 1;
  ram[11155]  = 1;
  ram[11156]  = 1;
  ram[11157]  = 1;
  ram[11158]  = 1;
  ram[11159]  = 1;
  ram[11160]  = 1;
  ram[11161]  = 1;
  ram[11162]  = 1;
  ram[11163]  = 1;
  ram[11164]  = 1;
  ram[11165]  = 1;
  ram[11166]  = 1;
  ram[11167]  = 1;
  ram[11168]  = 1;
  ram[11169]  = 1;
  ram[11170]  = 1;
  ram[11171]  = 1;
  ram[11172]  = 1;
  ram[11173]  = 1;
  ram[11174]  = 1;
  ram[11175]  = 1;
  ram[11176]  = 1;
  ram[11177]  = 1;
  ram[11178]  = 1;
  ram[11179]  = 1;
  ram[11180]  = 1;
  ram[11181]  = 1;
  ram[11182]  = 1;
  ram[11183]  = 1;
  ram[11184]  = 1;
  ram[11185]  = 1;
  ram[11186]  = 1;
  ram[11187]  = 1;
  ram[11188]  = 1;
  ram[11189]  = 1;
  ram[11190]  = 1;
  ram[11191]  = 1;
  ram[11192]  = 1;
  ram[11193]  = 1;
  ram[11194]  = 1;
  ram[11195]  = 1;
  ram[11196]  = 1;
  ram[11197]  = 1;
  ram[11198]  = 1;
  ram[11199]  = 1;
  ram[11200]  = 1;
  ram[11201]  = 1;
  ram[11202]  = 0;
  ram[11203]  = 0;
  ram[11204]  = 0;
  ram[11205]  = 1;
  ram[11206]  = 1;
  ram[11207]  = 0;
  ram[11208]  = 0;
  ram[11209]  = 1;
  ram[11210]  = 1;
  ram[11211]  = 1;
  ram[11212]  = 1;
  ram[11213]  = 0;
  ram[11214]  = 1;
  ram[11215]  = 1;
  ram[11216]  = 1;
  ram[11217]  = 0;
  ram[11218]  = 0;
  ram[11219]  = 1;
  ram[11220]  = 1;
  ram[11221]  = 1;
  ram[11222]  = 0;
  ram[11223]  = 0;
  ram[11224]  = 1;
  ram[11225]  = 1;
  ram[11226]  = 1;
  ram[11227]  = 1;
  ram[11228]  = 0;
  ram[11229]  = 1;
  ram[11230]  = 1;
  ram[11231]  = 1;
  ram[11232]  = 1;
  ram[11233]  = 1;
  ram[11234]  = 0;
  ram[11235]  = 1;
  ram[11236]  = 1;
  ram[11237]  = 1;
  ram[11238]  = 0;
  ram[11239]  = 0;
  ram[11240]  = 1;
  ram[11241]  = 1;
  ram[11242]  = 1;
  ram[11243]  = 0;
  ram[11244]  = 1;
  ram[11245]  = 1;
  ram[11246]  = 1;
  ram[11247]  = 1;
  ram[11248]  = 1;
  ram[11249]  = 1;
  ram[11250]  = 1;
  ram[11251]  = 1;
  ram[11252]  = 1;
  ram[11253]  = 1;
  ram[11254]  = 0;
  ram[11255]  = 0;
  ram[11256]  = 0;
  ram[11257]  = 1;
  ram[11258]  = 1;
  ram[11259]  = 0;
  ram[11260]  = 0;
  ram[11261]  = 0;
  ram[11262]  = 1;
  ram[11263]  = 1;
  ram[11264]  = 1;
  ram[11265]  = 1;
  ram[11266]  = 1;
  ram[11267]  = 1;
  ram[11268]  = 0;
  ram[11269]  = 0;
  ram[11270]  = 1;
  ram[11271]  = 1;
  ram[11272]  = 1;
  ram[11273]  = 1;
  ram[11274]  = 1;
  ram[11275]  = 1;
  ram[11276]  = 0;
  ram[11277]  = 0;
  ram[11278]  = 1;
  ram[11279]  = 1;
  ram[11280]  = 0;
  ram[11281]  = 0;
  ram[11282]  = 1;
  ram[11283]  = 1;
  ram[11284]  = 1;
  ram[11285]  = 0;
  ram[11286]  = 1;
  ram[11287]  = 1;
  ram[11288]  = 1;
  ram[11289]  = 1;
  ram[11290]  = 1;
  ram[11291]  = 0;
  ram[11292]  = 0;
  ram[11293]  = 1;
  ram[11294]  = 1;
  ram[11295]  = 1;
  ram[11296]  = 1;
  ram[11297]  = 1;
  ram[11298]  = 1;
  ram[11299]  = 1;
  ram[11300]  = 1;
  ram[11301]  = 1;
  ram[11302]  = 1;
  ram[11303]  = 1;
  ram[11304]  = 1;
  ram[11305]  = 1;
  ram[11306]  = 1;
  ram[11307]  = 1;
  ram[11308]  = 1;
  ram[11309]  = 1;
  ram[11310]  = 1;
  ram[11311]  = 1;
  ram[11312]  = 1;
  ram[11313]  = 1;
  ram[11314]  = 1;
  ram[11315]  = 1;
  ram[11316]  = 1;
  ram[11317]  = 1;
  ram[11318]  = 1;
  ram[11319]  = 1;
  ram[11320]  = 1;
  ram[11321]  = 1;
  ram[11322]  = 1;
  ram[11323]  = 1;
  ram[11324]  = 1;
  ram[11325]  = 1;
  ram[11326]  = 1;
  ram[11327]  = 1;
  ram[11328]  = 1;
  ram[11329]  = 1;
  ram[11330]  = 1;
  ram[11331]  = 1;
  ram[11332]  = 1;
  ram[11333]  = 1;
  ram[11334]  = 1;
  ram[11335]  = 1;
  ram[11336]  = 1;
  ram[11337]  = 1;
  ram[11338]  = 1;
  ram[11339]  = 1;
  ram[11340]  = 1;
  ram[11341]  = 1;
  ram[11342]  = 1;
  ram[11343]  = 1;
  ram[11344]  = 1;
  ram[11345]  = 1;
  ram[11346]  = 1;
  ram[11347]  = 1;
  ram[11348]  = 1;
  ram[11349]  = 1;
  ram[11350]  = 1;
  ram[11351]  = 1;
  ram[11352]  = 1;
  ram[11353]  = 1;
  ram[11354]  = 1;
  ram[11355]  = 1;
  ram[11356]  = 1;
  ram[11357]  = 1;
  ram[11358]  = 1;
  ram[11359]  = 1;
  ram[11360]  = 1;
  ram[11361]  = 1;
  ram[11362]  = 1;
  ram[11363]  = 1;
  ram[11364]  = 1;
  ram[11365]  = 1;
  ram[11366]  = 1;
  ram[11367]  = 1;
  ram[11368]  = 1;
  ram[11369]  = 1;
  ram[11370]  = 1;
  ram[11371]  = 1;
  ram[11372]  = 1;
  ram[11373]  = 1;
  ram[11374]  = 1;
  ram[11375]  = 1;
  ram[11376]  = 1;
  ram[11377]  = 1;
  ram[11378]  = 1;
  ram[11379]  = 1;
  ram[11380]  = 1;
  ram[11381]  = 1;
  ram[11382]  = 1;
  ram[11383]  = 1;
  ram[11384]  = 1;
  ram[11385]  = 1;
  ram[11386]  = 1;
  ram[11387]  = 1;
  ram[11388]  = 1;
  ram[11389]  = 1;
  ram[11390]  = 1;
  ram[11391]  = 1;
  ram[11392]  = 1;
  ram[11393]  = 1;
  ram[11394]  = 1;
  ram[11395]  = 1;
  ram[11396]  = 1;
  ram[11397]  = 1;
  ram[11398]  = 1;
  ram[11399]  = 1;
  ram[11400]  = 1;
  ram[11401]  = 1;
  ram[11402]  = 1;
  ram[11403]  = 1;
  ram[11404]  = 1;
  ram[11405]  = 1;
  ram[11406]  = 1;
  ram[11407]  = 1;
  ram[11408]  = 1;
  ram[11409]  = 1;
  ram[11410]  = 1;
  ram[11411]  = 1;
  ram[11412]  = 1;
  ram[11413]  = 1;
  ram[11414]  = 1;
  ram[11415]  = 1;
  ram[11416]  = 1;
  ram[11417]  = 1;
  ram[11418]  = 1;
  ram[11419]  = 1;
  ram[11420]  = 1;
  ram[11421]  = 1;
  ram[11422]  = 1;
  ram[11423]  = 1;
  ram[11424]  = 1;
  ram[11425]  = 1;
  ram[11426]  = 1;
  ram[11427]  = 1;
  ram[11428]  = 1;
  ram[11429]  = 1;
  ram[11430]  = 1;
  ram[11431]  = 1;
  ram[11432]  = 1;
  ram[11433]  = 1;
  ram[11434]  = 1;
  ram[11435]  = 1;
  ram[11436]  = 1;
  ram[11437]  = 1;
  ram[11438]  = 1;
  ram[11439]  = 1;
  ram[11440]  = 1;
  ram[11441]  = 1;
  ram[11442]  = 1;
  ram[11443]  = 1;
  ram[11444]  = 1;
  ram[11445]  = 1;
  ram[11446]  = 1;
  ram[11447]  = 1;
  ram[11448]  = 1;
  ram[11449]  = 1;
  ram[11450]  = 1;
  ram[11451]  = 1;
  ram[11452]  = 1;
  ram[11453]  = 1;
  ram[11454]  = 1;
  ram[11455]  = 1;
  ram[11456]  = 1;
  ram[11457]  = 1;
  ram[11458]  = 1;
  ram[11459]  = 1;
  ram[11460]  = 1;
  ram[11461]  = 1;
  ram[11462]  = 1;
  ram[11463]  = 1;
  ram[11464]  = 1;
  ram[11465]  = 1;
  ram[11466]  = 1;
  ram[11467]  = 1;
  ram[11468]  = 1;
  ram[11469]  = 1;
  ram[11470]  = 1;
  ram[11471]  = 1;
  ram[11472]  = 1;
  ram[11473]  = 1;
  ram[11474]  = 1;
  ram[11475]  = 1;
  ram[11476]  = 1;
  ram[11477]  = 1;
  ram[11478]  = 1;
  ram[11479]  = 1;
  ram[11480]  = 1;
  ram[11481]  = 1;
  ram[11482]  = 1;
  ram[11483]  = 1;
  ram[11484]  = 1;
  ram[11485]  = 1;
  ram[11486]  = 1;
  ram[11487]  = 1;
  ram[11488]  = 1;
  ram[11489]  = 1;
  ram[11490]  = 1;
  ram[11491]  = 1;
  ram[11492]  = 1;
  ram[11493]  = 1;
  ram[11494]  = 1;
  ram[11495]  = 1;
  ram[11496]  = 1;
  ram[11497]  = 1;
  ram[11498]  = 1;
  ram[11499]  = 1;
  ram[11500]  = 1;
  ram[11501]  = 1;
  ram[11502]  = 1;
  ram[11503]  = 0;
  ram[11504]  = 0;
  ram[11505]  = 0;
  ram[11506]  = 0;
  ram[11507]  = 0;
  ram[11508]  = 1;
  ram[11509]  = 1;
  ram[11510]  = 1;
  ram[11511]  = 1;
  ram[11512]  = 1;
  ram[11513]  = 0;
  ram[11514]  = 0;
  ram[11515]  = 0;
  ram[11516]  = 0;
  ram[11517]  = 1;
  ram[11518]  = 0;
  ram[11519]  = 0;
  ram[11520]  = 1;
  ram[11521]  = 1;
  ram[11522]  = 0;
  ram[11523]  = 0;
  ram[11524]  = 1;
  ram[11525]  = 1;
  ram[11526]  = 1;
  ram[11527]  = 1;
  ram[11528]  = 0;
  ram[11529]  = 1;
  ram[11530]  = 1;
  ram[11531]  = 1;
  ram[11532]  = 1;
  ram[11533]  = 1;
  ram[11534]  = 0;
  ram[11535]  = 1;
  ram[11536]  = 1;
  ram[11537]  = 1;
  ram[11538]  = 1;
  ram[11539]  = 0;
  ram[11540]  = 0;
  ram[11541]  = 0;
  ram[11542]  = 0;
  ram[11543]  = 0;
  ram[11544]  = 1;
  ram[11545]  = 1;
  ram[11546]  = 1;
  ram[11547]  = 1;
  ram[11548]  = 1;
  ram[11549]  = 1;
  ram[11550]  = 1;
  ram[11551]  = 1;
  ram[11552]  = 1;
  ram[11553]  = 1;
  ram[11554]  = 1;
  ram[11555]  = 0;
  ram[11556]  = 0;
  ram[11557]  = 0;
  ram[11558]  = 0;
  ram[11559]  = 0;
  ram[11560]  = 0;
  ram[11561]  = 1;
  ram[11562]  = 1;
  ram[11563]  = 1;
  ram[11564]  = 1;
  ram[11565]  = 1;
  ram[11566]  = 1;
  ram[11567]  = 1;
  ram[11568]  = 0;
  ram[11569]  = 0;
  ram[11570]  = 1;
  ram[11571]  = 1;
  ram[11572]  = 1;
  ram[11573]  = 1;
  ram[11574]  = 1;
  ram[11575]  = 1;
  ram[11576]  = 0;
  ram[11577]  = 0;
  ram[11578]  = 0;
  ram[11579]  = 0;
  ram[11580]  = 0;
  ram[11581]  = 1;
  ram[11582]  = 1;
  ram[11583]  = 1;
  ram[11584]  = 1;
  ram[11585]  = 0;
  ram[11586]  = 1;
  ram[11587]  = 1;
  ram[11588]  = 1;
  ram[11589]  = 1;
  ram[11590]  = 1;
  ram[11591]  = 0;
  ram[11592]  = 0;
  ram[11593]  = 1;
  ram[11594]  = 1;
  ram[11595]  = 1;
  ram[11596]  = 1;
  ram[11597]  = 1;
  ram[11598]  = 1;
  ram[11599]  = 1;
  ram[11600]  = 1;
  ram[11601]  = 1;
  ram[11602]  = 1;
  ram[11603]  = 1;
  ram[11604]  = 1;
  ram[11605]  = 1;
  ram[11606]  = 1;
  ram[11607]  = 1;
  ram[11608]  = 1;
  ram[11609]  = 1;
  ram[11610]  = 1;
  ram[11611]  = 1;
  ram[11612]  = 1;
  ram[11613]  = 1;
  ram[11614]  = 1;
  ram[11615]  = 1;
  ram[11616]  = 1;
  ram[11617]  = 1;
  ram[11618]  = 1;
  ram[11619]  = 1;
  ram[11620]  = 1;
  ram[11621]  = 1;
  ram[11622]  = 1;
  ram[11623]  = 1;
  ram[11624]  = 1;
  ram[11625]  = 1;
  ram[11626]  = 1;
  ram[11627]  = 1;
  ram[11628]  = 1;
  ram[11629]  = 1;
  ram[11630]  = 1;
  ram[11631]  = 1;
  ram[11632]  = 1;
  ram[11633]  = 1;
  ram[11634]  = 1;
  ram[11635]  = 1;
  ram[11636]  = 1;
  ram[11637]  = 1;
  ram[11638]  = 1;
  ram[11639]  = 1;
  ram[11640]  = 1;
  ram[11641]  = 1;
  ram[11642]  = 1;
  ram[11643]  = 1;
  ram[11644]  = 1;
  ram[11645]  = 1;
  ram[11646]  = 1;
  ram[11647]  = 1;
  ram[11648]  = 1;
  ram[11649]  = 1;
  ram[11650]  = 1;
  ram[11651]  = 1;
  ram[11652]  = 1;
  ram[11653]  = 1;
  ram[11654]  = 1;
  ram[11655]  = 1;
  ram[11656]  = 1;
  ram[11657]  = 1;
  ram[11658]  = 1;
  ram[11659]  = 1;
  ram[11660]  = 1;
  ram[11661]  = 1;
  ram[11662]  = 1;
  ram[11663]  = 1;
  ram[11664]  = 1;
  ram[11665]  = 1;
  ram[11666]  = 1;
  ram[11667]  = 1;
  ram[11668]  = 1;
  ram[11669]  = 1;
  ram[11670]  = 1;
  ram[11671]  = 1;
  ram[11672]  = 1;
  ram[11673]  = 1;
  ram[11674]  = 1;
  ram[11675]  = 1;
  ram[11676]  = 1;
  ram[11677]  = 1;
  ram[11678]  = 1;
  ram[11679]  = 1;
  ram[11680]  = 1;
  ram[11681]  = 1;
  ram[11682]  = 1;
  ram[11683]  = 1;
  ram[11684]  = 1;
  ram[11685]  = 1;
  ram[11686]  = 1;
  ram[11687]  = 1;
  ram[11688]  = 1;
  ram[11689]  = 1;
  ram[11690]  = 1;
  ram[11691]  = 1;
  ram[11692]  = 1;
  ram[11693]  = 1;
  ram[11694]  = 1;
  ram[11695]  = 1;
  ram[11696]  = 1;
  ram[11697]  = 1;
  ram[11698]  = 1;
  ram[11699]  = 1;
  ram[11700]  = 1;
  ram[11701]  = 1;
  ram[11702]  = 1;
  ram[11703]  = 1;
  ram[11704]  = 1;
  ram[11705]  = 1;
  ram[11706]  = 1;
  ram[11707]  = 1;
  ram[11708]  = 1;
  ram[11709]  = 1;
  ram[11710]  = 1;
  ram[11711]  = 1;
  ram[11712]  = 1;
  ram[11713]  = 1;
  ram[11714]  = 1;
  ram[11715]  = 1;
  ram[11716]  = 1;
  ram[11717]  = 1;
  ram[11718]  = 1;
  ram[11719]  = 1;
  ram[11720]  = 1;
  ram[11721]  = 1;
  ram[11722]  = 1;
  ram[11723]  = 1;
  ram[11724]  = 1;
  ram[11725]  = 1;
  ram[11726]  = 1;
  ram[11727]  = 1;
  ram[11728]  = 1;
  ram[11729]  = 1;
  ram[11730]  = 1;
  ram[11731]  = 1;
  ram[11732]  = 1;
  ram[11733]  = 1;
  ram[11734]  = 1;
  ram[11735]  = 1;
  ram[11736]  = 1;
  ram[11737]  = 1;
  ram[11738]  = 1;
  ram[11739]  = 1;
  ram[11740]  = 1;
  ram[11741]  = 1;
  ram[11742]  = 1;
  ram[11743]  = 1;
  ram[11744]  = 1;
  ram[11745]  = 1;
  ram[11746]  = 1;
  ram[11747]  = 1;
  ram[11748]  = 1;
  ram[11749]  = 1;
  ram[11750]  = 1;
  ram[11751]  = 1;
  ram[11752]  = 1;
  ram[11753]  = 1;
  ram[11754]  = 1;
  ram[11755]  = 1;
  ram[11756]  = 1;
  ram[11757]  = 1;
  ram[11758]  = 1;
  ram[11759]  = 1;
  ram[11760]  = 1;
  ram[11761]  = 1;
  ram[11762]  = 1;
  ram[11763]  = 1;
  ram[11764]  = 1;
  ram[11765]  = 1;
  ram[11766]  = 1;
  ram[11767]  = 1;
  ram[11768]  = 1;
  ram[11769]  = 1;
  ram[11770]  = 1;
  ram[11771]  = 1;
  ram[11772]  = 1;
  ram[11773]  = 1;
  ram[11774]  = 1;
  ram[11775]  = 1;
  ram[11776]  = 1;
  ram[11777]  = 1;
  ram[11778]  = 1;
  ram[11779]  = 1;
  ram[11780]  = 1;
  ram[11781]  = 1;
  ram[11782]  = 1;
  ram[11783]  = 1;
  ram[11784]  = 1;
  ram[11785]  = 1;
  ram[11786]  = 1;
  ram[11787]  = 1;
  ram[11788]  = 1;
  ram[11789]  = 1;
  ram[11790]  = 1;
  ram[11791]  = 1;
  ram[11792]  = 1;
  ram[11793]  = 1;
  ram[11794]  = 1;
  ram[11795]  = 1;
  ram[11796]  = 1;
  ram[11797]  = 1;
  ram[11798]  = 1;
  ram[11799]  = 1;
  ram[11800]  = 1;
  ram[11801]  = 1;
  ram[11802]  = 1;
  ram[11803]  = 1;
  ram[11804]  = 1;
  ram[11805]  = 0;
  ram[11806]  = 1;
  ram[11807]  = 1;
  ram[11808]  = 1;
  ram[11809]  = 1;
  ram[11810]  = 1;
  ram[11811]  = 1;
  ram[11812]  = 1;
  ram[11813]  = 1;
  ram[11814]  = 1;
  ram[11815]  = 0;
  ram[11816]  = 1;
  ram[11817]  = 1;
  ram[11818]  = 1;
  ram[11819]  = 1;
  ram[11820]  = 1;
  ram[11821]  = 1;
  ram[11822]  = 1;
  ram[11823]  = 1;
  ram[11824]  = 1;
  ram[11825]  = 1;
  ram[11826]  = 1;
  ram[11827]  = 1;
  ram[11828]  = 1;
  ram[11829]  = 1;
  ram[11830]  = 1;
  ram[11831]  = 1;
  ram[11832]  = 1;
  ram[11833]  = 1;
  ram[11834]  = 1;
  ram[11835]  = 1;
  ram[11836]  = 1;
  ram[11837]  = 1;
  ram[11838]  = 1;
  ram[11839]  = 1;
  ram[11840]  = 1;
  ram[11841]  = 0;
  ram[11842]  = 1;
  ram[11843]  = 1;
  ram[11844]  = 1;
  ram[11845]  = 1;
  ram[11846]  = 1;
  ram[11847]  = 1;
  ram[11848]  = 1;
  ram[11849]  = 1;
  ram[11850]  = 1;
  ram[11851]  = 1;
  ram[11852]  = 1;
  ram[11853]  = 1;
  ram[11854]  = 1;
  ram[11855]  = 1;
  ram[11856]  = 1;
  ram[11857]  = 1;
  ram[11858]  = 0;
  ram[11859]  = 1;
  ram[11860]  = 1;
  ram[11861]  = 1;
  ram[11862]  = 1;
  ram[11863]  = 1;
  ram[11864]  = 1;
  ram[11865]  = 1;
  ram[11866]  = 1;
  ram[11867]  = 1;
  ram[11868]  = 1;
  ram[11869]  = 1;
  ram[11870]  = 1;
  ram[11871]  = 1;
  ram[11872]  = 1;
  ram[11873]  = 1;
  ram[11874]  = 1;
  ram[11875]  = 1;
  ram[11876]  = 1;
  ram[11877]  = 1;
  ram[11878]  = 0;
  ram[11879]  = 1;
  ram[11880]  = 1;
  ram[11881]  = 1;
  ram[11882]  = 1;
  ram[11883]  = 1;
  ram[11884]  = 1;
  ram[11885]  = 1;
  ram[11886]  = 1;
  ram[11887]  = 1;
  ram[11888]  = 1;
  ram[11889]  = 1;
  ram[11890]  = 1;
  ram[11891]  = 1;
  ram[11892]  = 1;
  ram[11893]  = 1;
  ram[11894]  = 1;
  ram[11895]  = 1;
  ram[11896]  = 1;
  ram[11897]  = 1;
  ram[11898]  = 1;
  ram[11899]  = 1;
  ram[11900]  = 1;
  ram[11901]  = 1;
  ram[11902]  = 1;
  ram[11903]  = 1;
  ram[11904]  = 1;
  ram[11905]  = 1;
  ram[11906]  = 1;
  ram[11907]  = 1;
  ram[11908]  = 1;
  ram[11909]  = 1;
  ram[11910]  = 1;
  ram[11911]  = 1;
  ram[11912]  = 1;
  ram[11913]  = 1;
  ram[11914]  = 1;
  ram[11915]  = 1;
  ram[11916]  = 1;
  ram[11917]  = 1;
  ram[11918]  = 1;
  ram[11919]  = 1;
  ram[11920]  = 1;
  ram[11921]  = 1;
  ram[11922]  = 1;
  ram[11923]  = 1;
  ram[11924]  = 1;
  ram[11925]  = 1;
  ram[11926]  = 1;
  ram[11927]  = 1;
  ram[11928]  = 1;
  ram[11929]  = 1;
  ram[11930]  = 1;
  ram[11931]  = 1;
  ram[11932]  = 1;
  ram[11933]  = 1;
  ram[11934]  = 1;
  ram[11935]  = 1;
  ram[11936]  = 1;
  ram[11937]  = 1;
  ram[11938]  = 1;
  ram[11939]  = 1;
  ram[11940]  = 1;
  ram[11941]  = 1;
  ram[11942]  = 1;
  ram[11943]  = 1;
  ram[11944]  = 1;
  ram[11945]  = 1;
  ram[11946]  = 1;
  ram[11947]  = 1;
  ram[11948]  = 1;
  ram[11949]  = 1;
  ram[11950]  = 1;
  ram[11951]  = 1;
  ram[11952]  = 1;
  ram[11953]  = 1;
  ram[11954]  = 1;
  ram[11955]  = 1;
  ram[11956]  = 1;
  ram[11957]  = 1;
  ram[11958]  = 1;
  ram[11959]  = 1;
  ram[11960]  = 1;
  ram[11961]  = 1;
  ram[11962]  = 1;
  ram[11963]  = 1;
  ram[11964]  = 1;
  ram[11965]  = 1;
  ram[11966]  = 1;
  ram[11967]  = 1;
  ram[11968]  = 1;
  ram[11969]  = 1;
  ram[11970]  = 1;
  ram[11971]  = 1;
  ram[11972]  = 1;
  ram[11973]  = 1;
  ram[11974]  = 1;
  ram[11975]  = 1;
  ram[11976]  = 1;
  ram[11977]  = 1;
  ram[11978]  = 1;
  ram[11979]  = 1;
  ram[11980]  = 1;
  ram[11981]  = 1;
  ram[11982]  = 1;
  ram[11983]  = 1;
  ram[11984]  = 1;
  ram[11985]  = 1;
  ram[11986]  = 1;
  ram[11987]  = 1;
  ram[11988]  = 1;
  ram[11989]  = 1;
  ram[11990]  = 1;
  ram[11991]  = 1;
  ram[11992]  = 1;
  ram[11993]  = 1;
  ram[11994]  = 1;
  ram[11995]  = 1;
  ram[11996]  = 1;
  ram[11997]  = 1;
  ram[11998]  = 1;
  ram[11999]  = 1;
  ram[12000]  = 1;
  ram[12001]  = 1;
  ram[12002]  = 1;
  ram[12003]  = 1;
  ram[12004]  = 1;
  ram[12005]  = 1;
  ram[12006]  = 1;
  ram[12007]  = 1;
  ram[12008]  = 1;
  ram[12009]  = 1;
  ram[12010]  = 1;
  ram[12011]  = 1;
  ram[12012]  = 1;
  ram[12013]  = 1;
  ram[12014]  = 1;
  ram[12015]  = 1;
  ram[12016]  = 1;
  ram[12017]  = 1;
  ram[12018]  = 1;
  ram[12019]  = 1;
  ram[12020]  = 1;
  ram[12021]  = 1;
  ram[12022]  = 1;
  ram[12023]  = 1;
  ram[12024]  = 1;
  ram[12025]  = 1;
  ram[12026]  = 1;
  ram[12027]  = 1;
  ram[12028]  = 1;
  ram[12029]  = 1;
  ram[12030]  = 1;
  ram[12031]  = 1;
  ram[12032]  = 1;
  ram[12033]  = 1;
  ram[12034]  = 1;
  ram[12035]  = 1;
  ram[12036]  = 1;
  ram[12037]  = 1;
  ram[12038]  = 1;
  ram[12039]  = 1;
  ram[12040]  = 1;
  ram[12041]  = 1;
  ram[12042]  = 1;
  ram[12043]  = 1;
  ram[12044]  = 1;
  ram[12045]  = 1;
  ram[12046]  = 1;
  ram[12047]  = 1;
  ram[12048]  = 1;
  ram[12049]  = 1;
  ram[12050]  = 1;
  ram[12051]  = 1;
  ram[12052]  = 1;
  ram[12053]  = 1;
  ram[12054]  = 1;
  ram[12055]  = 1;
  ram[12056]  = 1;
  ram[12057]  = 1;
  ram[12058]  = 1;
  ram[12059]  = 1;
  ram[12060]  = 1;
  ram[12061]  = 1;
  ram[12062]  = 1;
  ram[12063]  = 1;
  ram[12064]  = 1;
  ram[12065]  = 1;
  ram[12066]  = 1;
  ram[12067]  = 1;
  ram[12068]  = 1;
  ram[12069]  = 1;
  ram[12070]  = 1;
  ram[12071]  = 1;
  ram[12072]  = 1;
  ram[12073]  = 1;
  ram[12074]  = 1;
  ram[12075]  = 1;
  ram[12076]  = 1;
  ram[12077]  = 1;
  ram[12078]  = 1;
  ram[12079]  = 1;
  ram[12080]  = 1;
  ram[12081]  = 1;
  ram[12082]  = 1;
  ram[12083]  = 1;
  ram[12084]  = 1;
  ram[12085]  = 1;
  ram[12086]  = 1;
  ram[12087]  = 1;
  ram[12088]  = 1;
  ram[12089]  = 1;
  ram[12090]  = 1;
  ram[12091]  = 1;
  ram[12092]  = 1;
  ram[12093]  = 1;
  ram[12094]  = 1;
  ram[12095]  = 1;
  ram[12096]  = 1;
  ram[12097]  = 1;
  ram[12098]  = 1;
  ram[12099]  = 1;
  ram[12100]  = 1;
  ram[12101]  = 1;
  ram[12102]  = 1;
  ram[12103]  = 1;
  ram[12104]  = 1;
  ram[12105]  = 1;
  ram[12106]  = 1;
  ram[12107]  = 1;
  ram[12108]  = 1;
  ram[12109]  = 1;
  ram[12110]  = 1;
  ram[12111]  = 1;
  ram[12112]  = 1;
  ram[12113]  = 1;
  ram[12114]  = 1;
  ram[12115]  = 1;
  ram[12116]  = 1;
  ram[12117]  = 1;
  ram[12118]  = 1;
  ram[12119]  = 1;
  ram[12120]  = 1;
  ram[12121]  = 1;
  ram[12122]  = 1;
  ram[12123]  = 1;
  ram[12124]  = 1;
  ram[12125]  = 1;
  ram[12126]  = 1;
  ram[12127]  = 1;
  ram[12128]  = 1;
  ram[12129]  = 1;
  ram[12130]  = 1;
  ram[12131]  = 1;
  ram[12132]  = 1;
  ram[12133]  = 1;
  ram[12134]  = 1;
  ram[12135]  = 1;
  ram[12136]  = 1;
  ram[12137]  = 1;
  ram[12138]  = 1;
  ram[12139]  = 1;
  ram[12140]  = 1;
  ram[12141]  = 1;
  ram[12142]  = 1;
  ram[12143]  = 1;
  ram[12144]  = 1;
  ram[12145]  = 1;
  ram[12146]  = 1;
  ram[12147]  = 1;
  ram[12148]  = 1;
  ram[12149]  = 1;
  ram[12150]  = 1;
  ram[12151]  = 1;
  ram[12152]  = 1;
  ram[12153]  = 1;
  ram[12154]  = 1;
  ram[12155]  = 1;
  ram[12156]  = 1;
  ram[12157]  = 1;
  ram[12158]  = 1;
  ram[12159]  = 1;
  ram[12160]  = 1;
  ram[12161]  = 1;
  ram[12162]  = 1;
  ram[12163]  = 1;
  ram[12164]  = 1;
  ram[12165]  = 1;
  ram[12166]  = 1;
  ram[12167]  = 1;
  ram[12168]  = 1;
  ram[12169]  = 1;
  ram[12170]  = 1;
  ram[12171]  = 1;
  ram[12172]  = 1;
  ram[12173]  = 1;
  ram[12174]  = 1;
  ram[12175]  = 1;
  ram[12176]  = 1;
  ram[12177]  = 1;
  ram[12178]  = 1;
  ram[12179]  = 1;
  ram[12180]  = 1;
  ram[12181]  = 1;
  ram[12182]  = 1;
  ram[12183]  = 1;
  ram[12184]  = 1;
  ram[12185]  = 1;
  ram[12186]  = 1;
  ram[12187]  = 1;
  ram[12188]  = 1;
  ram[12189]  = 1;
  ram[12190]  = 1;
  ram[12191]  = 1;
  ram[12192]  = 1;
  ram[12193]  = 1;
  ram[12194]  = 1;
  ram[12195]  = 1;
  ram[12196]  = 1;
  ram[12197]  = 1;
  ram[12198]  = 1;
  ram[12199]  = 1;
  ram[12200]  = 1;
  ram[12201]  = 1;
  ram[12202]  = 1;
  ram[12203]  = 1;
  ram[12204]  = 1;
  ram[12205]  = 1;
  ram[12206]  = 1;
  ram[12207]  = 1;
  ram[12208]  = 1;
  ram[12209]  = 1;
  ram[12210]  = 1;
  ram[12211]  = 1;
  ram[12212]  = 1;
  ram[12213]  = 1;
  ram[12214]  = 1;
  ram[12215]  = 1;
  ram[12216]  = 1;
  ram[12217]  = 1;
  ram[12218]  = 1;
  ram[12219]  = 1;
  ram[12220]  = 1;
  ram[12221]  = 1;
  ram[12222]  = 1;
  ram[12223]  = 1;
  ram[12224]  = 1;
  ram[12225]  = 1;
  ram[12226]  = 1;
  ram[12227]  = 1;
  ram[12228]  = 1;
  ram[12229]  = 1;
  ram[12230]  = 1;
  ram[12231]  = 1;
  ram[12232]  = 1;
  ram[12233]  = 1;
  ram[12234]  = 1;
  ram[12235]  = 1;
  ram[12236]  = 1;
  ram[12237]  = 1;
  ram[12238]  = 1;
  ram[12239]  = 1;
  ram[12240]  = 1;
  ram[12241]  = 1;
  ram[12242]  = 1;
  ram[12243]  = 1;
  ram[12244]  = 1;
  ram[12245]  = 1;
  ram[12246]  = 1;
  ram[12247]  = 1;
  ram[12248]  = 1;
  ram[12249]  = 1;
  ram[12250]  = 1;
  ram[12251]  = 1;
  ram[12252]  = 1;
  ram[12253]  = 1;
  ram[12254]  = 1;
  ram[12255]  = 1;
  ram[12256]  = 1;
  ram[12257]  = 1;
  ram[12258]  = 1;
  ram[12259]  = 1;
  ram[12260]  = 1;
  ram[12261]  = 1;
  ram[12262]  = 1;
  ram[12263]  = 1;
  ram[12264]  = 1;
  ram[12265]  = 1;
  ram[12266]  = 1;
  ram[12267]  = 1;
  ram[12268]  = 1;
  ram[12269]  = 1;
  ram[12270]  = 1;
  ram[12271]  = 1;
  ram[12272]  = 1;
  ram[12273]  = 1;
  ram[12274]  = 1;
  ram[12275]  = 1;
  ram[12276]  = 1;
  ram[12277]  = 1;
  ram[12278]  = 1;
  ram[12279]  = 1;
  ram[12280]  = 1;
  ram[12281]  = 1;
  ram[12282]  = 1;
  ram[12283]  = 1;
  ram[12284]  = 1;
  ram[12285]  = 1;
  ram[12286]  = 1;
  ram[12287]  = 1;
  ram[12288]  = 1;
  ram[12289]  = 1;
  ram[12290]  = 1;
  ram[12291]  = 1;
  ram[12292]  = 1;
  ram[12293]  = 1;
  ram[12294]  = 1;
  ram[12295]  = 1;
  ram[12296]  = 1;
  ram[12297]  = 1;
  ram[12298]  = 1;
  ram[12299]  = 1;
  ram[12300]  = 1;
  ram[12301]  = 1;
  ram[12302]  = 1;
  ram[12303]  = 1;
  ram[12304]  = 1;
  ram[12305]  = 1;
  ram[12306]  = 1;
  ram[12307]  = 1;
  ram[12308]  = 1;
  ram[12309]  = 1;
  ram[12310]  = 1;
  ram[12311]  = 1;
  ram[12312]  = 1;
  ram[12313]  = 1;
  ram[12314]  = 1;
  ram[12315]  = 1;
  ram[12316]  = 1;
  ram[12317]  = 1;
  ram[12318]  = 1;
  ram[12319]  = 1;
  ram[12320]  = 1;
  ram[12321]  = 1;
  ram[12322]  = 1;
  ram[12323]  = 1;
  ram[12324]  = 1;
  ram[12325]  = 1;
  ram[12326]  = 1;
  ram[12327]  = 1;
  ram[12328]  = 1;
  ram[12329]  = 1;
  ram[12330]  = 1;
  ram[12331]  = 1;
  ram[12332]  = 1;
  ram[12333]  = 1;
  ram[12334]  = 1;
  ram[12335]  = 1;
  ram[12336]  = 1;
  ram[12337]  = 1;
  ram[12338]  = 1;
  ram[12339]  = 1;
  ram[12340]  = 1;
  ram[12341]  = 1;
  ram[12342]  = 1;
  ram[12343]  = 1;
  ram[12344]  = 1;
  ram[12345]  = 1;
  ram[12346]  = 1;
  ram[12347]  = 1;
  ram[12348]  = 1;
  ram[12349]  = 1;
  ram[12350]  = 1;
  ram[12351]  = 1;
  ram[12352]  = 1;
  ram[12353]  = 1;
  ram[12354]  = 1;
  ram[12355]  = 1;
  ram[12356]  = 1;
  ram[12357]  = 1;
  ram[12358]  = 1;
  ram[12359]  = 1;
  ram[12360]  = 1;
  ram[12361]  = 1;
  ram[12362]  = 1;
  ram[12363]  = 1;
  ram[12364]  = 1;
  ram[12365]  = 1;
  ram[12366]  = 1;
  ram[12367]  = 1;
  ram[12368]  = 1;
  ram[12369]  = 1;
  ram[12370]  = 1;
  ram[12371]  = 1;
  ram[12372]  = 1;
  ram[12373]  = 1;
  ram[12374]  = 1;
  ram[12375]  = 1;
  ram[12376]  = 1;
  ram[12377]  = 1;
  ram[12378]  = 1;
  ram[12379]  = 1;
  ram[12380]  = 1;
  ram[12381]  = 1;
  ram[12382]  = 1;
  ram[12383]  = 1;
  ram[12384]  = 1;
  ram[12385]  = 1;
  ram[12386]  = 1;
  ram[12387]  = 1;
  ram[12388]  = 1;
  ram[12389]  = 1;
  ram[12390]  = 1;
  ram[12391]  = 1;
  ram[12392]  = 1;
  ram[12393]  = 1;
  ram[12394]  = 1;
  ram[12395]  = 1;
  ram[12396]  = 1;
  ram[12397]  = 1;
  ram[12398]  = 1;
  ram[12399]  = 1;
  ram[12400]  = 1;
  ram[12401]  = 1;
  ram[12402]  = 1;
  ram[12403]  = 1;
  ram[12404]  = 1;
  ram[12405]  = 1;
  ram[12406]  = 1;
  ram[12407]  = 1;
  ram[12408]  = 1;
  ram[12409]  = 1;
  ram[12410]  = 1;
  ram[12411]  = 1;
  ram[12412]  = 1;
  ram[12413]  = 1;
  ram[12414]  = 1;
  ram[12415]  = 1;
  ram[12416]  = 1;
  ram[12417]  = 1;
  ram[12418]  = 1;
  ram[12419]  = 1;
  ram[12420]  = 1;
  ram[12421]  = 1;
  ram[12422]  = 1;
  ram[12423]  = 1;
  ram[12424]  = 1;
  ram[12425]  = 1;
  ram[12426]  = 1;
  ram[12427]  = 1;
  ram[12428]  = 1;
  ram[12429]  = 1;
  ram[12430]  = 1;
  ram[12431]  = 1;
  ram[12432]  = 1;
  ram[12433]  = 1;
  ram[12434]  = 1;
  ram[12435]  = 1;
  ram[12436]  = 1;
  ram[12437]  = 1;
  ram[12438]  = 1;
  ram[12439]  = 1;
  ram[12440]  = 1;
  ram[12441]  = 1;
  ram[12442]  = 1;
  ram[12443]  = 1;
  ram[12444]  = 1;
  ram[12445]  = 1;
  ram[12446]  = 1;
  ram[12447]  = 1;
  ram[12448]  = 1;
  ram[12449]  = 1;
  ram[12450]  = 1;
  ram[12451]  = 1;
  ram[12452]  = 1;
  ram[12453]  = 1;
  ram[12454]  = 1;
  ram[12455]  = 1;
  ram[12456]  = 1;
  ram[12457]  = 1;
  ram[12458]  = 1;
  ram[12459]  = 1;
  ram[12460]  = 1;
  ram[12461]  = 1;
  ram[12462]  = 1;
  ram[12463]  = 1;
  ram[12464]  = 1;
  ram[12465]  = 1;
  ram[12466]  = 1;
  ram[12467]  = 1;
  ram[12468]  = 1;
  ram[12469]  = 1;
  ram[12470]  = 1;
  ram[12471]  = 1;
  ram[12472]  = 1;
  ram[12473]  = 1;
  ram[12474]  = 1;
  ram[12475]  = 1;
  ram[12476]  = 1;
  ram[12477]  = 1;
  ram[12478]  = 1;
  ram[12479]  = 1;
  ram[12480]  = 1;
  ram[12481]  = 1;
  ram[12482]  = 1;
  ram[12483]  = 1;
  ram[12484]  = 1;
  ram[12485]  = 1;
  ram[12486]  = 1;
  ram[12487]  = 1;
  ram[12488]  = 1;
  ram[12489]  = 1;
  ram[12490]  = 1;
  ram[12491]  = 1;
  ram[12492]  = 1;
  ram[12493]  = 1;
  ram[12494]  = 1;
  ram[12495]  = 1;
  ram[12496]  = 1;
  ram[12497]  = 1;
  ram[12498]  = 1;
  ram[12499]  = 1;
  ram[12500]  = 1;
  ram[12501]  = 1;
  ram[12502]  = 1;
  ram[12503]  = 1;
  ram[12504]  = 1;
  ram[12505]  = 1;
  ram[12506]  = 1;
  ram[12507]  = 1;
  ram[12508]  = 1;
  ram[12509]  = 1;
  ram[12510]  = 1;
  ram[12511]  = 1;
  ram[12512]  = 1;
  ram[12513]  = 1;
  ram[12514]  = 1;
  ram[12515]  = 1;
  ram[12516]  = 1;
  ram[12517]  = 1;
  ram[12518]  = 1;
  ram[12519]  = 1;
  ram[12520]  = 1;
  ram[12521]  = 1;
  ram[12522]  = 1;
  ram[12523]  = 1;
  ram[12524]  = 1;
  ram[12525]  = 1;
  ram[12526]  = 1;
  ram[12527]  = 1;
  ram[12528]  = 1;
  ram[12529]  = 1;
  ram[12530]  = 1;
  ram[12531]  = 1;
  ram[12532]  = 1;
  ram[12533]  = 1;
  ram[12534]  = 1;
  ram[12535]  = 1;
  ram[12536]  = 1;
  ram[12537]  = 1;
  ram[12538]  = 1;
  ram[12539]  = 1;
  ram[12540]  = 1;
  ram[12541]  = 1;
  ram[12542]  = 1;
  ram[12543]  = 1;
  ram[12544]  = 1;
  ram[12545]  = 1;
  ram[12546]  = 1;
  ram[12547]  = 1;
  ram[12548]  = 1;
  ram[12549]  = 1;
  ram[12550]  = 1;
  ram[12551]  = 1;
  ram[12552]  = 1;
  ram[12553]  = 1;
  ram[12554]  = 1;
  ram[12555]  = 1;
  ram[12556]  = 1;
  ram[12557]  = 1;
  ram[12558]  = 1;
  ram[12559]  = 1;
  ram[12560]  = 1;
  ram[12561]  = 1;
  ram[12562]  = 1;
  ram[12563]  = 1;
  ram[12564]  = 1;
  ram[12565]  = 1;
  ram[12566]  = 1;
  ram[12567]  = 1;
  ram[12568]  = 1;
  ram[12569]  = 1;
  ram[12570]  = 1;
  ram[12571]  = 1;
  ram[12572]  = 1;
  ram[12573]  = 1;
  ram[12574]  = 1;
  ram[12575]  = 1;
  ram[12576]  = 1;
  ram[12577]  = 1;
  ram[12578]  = 1;
  ram[12579]  = 1;
  ram[12580]  = 1;
  ram[12581]  = 1;
  ram[12582]  = 1;
  ram[12583]  = 1;
  ram[12584]  = 1;
  ram[12585]  = 1;
  ram[12586]  = 1;
  ram[12587]  = 1;
  ram[12588]  = 1;
  ram[12589]  = 1;
  ram[12590]  = 1;
  ram[12591]  = 1;
  ram[12592]  = 1;
  ram[12593]  = 1;
  ram[12594]  = 1;
  ram[12595]  = 1;
  ram[12596]  = 1;
  ram[12597]  = 1;
  ram[12598]  = 1;
  ram[12599]  = 1;
  ram[12600]  = 1;
  ram[12601]  = 1;
  ram[12602]  = 1;
  ram[12603]  = 1;
  ram[12604]  = 1;
  ram[12605]  = 1;
  ram[12606]  = 1;
  ram[12607]  = 1;
  ram[12608]  = 1;
  ram[12609]  = 1;
  ram[12610]  = 1;
  ram[12611]  = 1;
  ram[12612]  = 1;
  ram[12613]  = 1;
  ram[12614]  = 1;
  ram[12615]  = 1;
  ram[12616]  = 1;
  ram[12617]  = 1;
  ram[12618]  = 1;
  ram[12619]  = 1;
  ram[12620]  = 1;
  ram[12621]  = 1;
  ram[12622]  = 1;
  ram[12623]  = 1;
  ram[12624]  = 1;
  ram[12625]  = 1;
  ram[12626]  = 1;
  ram[12627]  = 1;
  ram[12628]  = 1;
  ram[12629]  = 1;
  ram[12630]  = 1;
  ram[12631]  = 1;
  ram[12632]  = 1;
  ram[12633]  = 1;
  ram[12634]  = 1;
  ram[12635]  = 1;
  ram[12636]  = 1;
  ram[12637]  = 1;
  ram[12638]  = 1;
  ram[12639]  = 1;
  ram[12640]  = 1;
  ram[12641]  = 1;
  ram[12642]  = 1;
  ram[12643]  = 1;
  ram[12644]  = 1;
  ram[12645]  = 1;
  ram[12646]  = 1;
  ram[12647]  = 1;
  ram[12648]  = 1;
  ram[12649]  = 1;
  ram[12650]  = 1;
  ram[12651]  = 1;
  ram[12652]  = 1;
  ram[12653]  = 1;
  ram[12654]  = 1;
  ram[12655]  = 1;
  ram[12656]  = 1;
  ram[12657]  = 1;
  ram[12658]  = 1;
  ram[12659]  = 1;
  ram[12660]  = 1;
  ram[12661]  = 1;
  ram[12662]  = 1;
  ram[12663]  = 1;
  ram[12664]  = 1;
  ram[12665]  = 1;
  ram[12666]  = 1;
  ram[12667]  = 1;
  ram[12668]  = 1;
  ram[12669]  = 1;
  ram[12670]  = 1;
  ram[12671]  = 1;
  ram[12672]  = 1;
  ram[12673]  = 1;
  ram[12674]  = 1;
  ram[12675]  = 1;
  ram[12676]  = 1;
  ram[12677]  = 1;
  ram[12678]  = 1;
  ram[12679]  = 1;
  ram[12680]  = 1;
  ram[12681]  = 1;
  ram[12682]  = 1;
  ram[12683]  = 1;
  ram[12684]  = 1;
  ram[12685]  = 1;
  ram[12686]  = 1;
  ram[12687]  = 1;
  ram[12688]  = 1;
  ram[12689]  = 1;
  ram[12690]  = 1;
  ram[12691]  = 1;
  ram[12692]  = 1;
  ram[12693]  = 1;
  ram[12694]  = 1;
  ram[12695]  = 1;
  ram[12696]  = 1;
  ram[12697]  = 1;
  ram[12698]  = 1;
  ram[12699]  = 1;
  ram[12700]  = 1;
  ram[12701]  = 1;
  ram[12702]  = 1;
  ram[12703]  = 1;
  ram[12704]  = 1;
  ram[12705]  = 1;
  ram[12706]  = 1;
  ram[12707]  = 1;
  ram[12708]  = 1;
  ram[12709]  = 1;
  ram[12710]  = 1;
  ram[12711]  = 1;
  ram[12712]  = 1;
  ram[12713]  = 1;
  ram[12714]  = 1;
  ram[12715]  = 1;
  ram[12716]  = 1;
  ram[12717]  = 1;
  ram[12718]  = 1;
  ram[12719]  = 1;
  ram[12720]  = 1;
  ram[12721]  = 1;
  ram[12722]  = 1;
  ram[12723]  = 1;
  ram[12724]  = 1;
  ram[12725]  = 1;
  ram[12726]  = 1;
  ram[12727]  = 1;
  ram[12728]  = 1;
  ram[12729]  = 1;
  ram[12730]  = 1;
  ram[12731]  = 1;
  ram[12732]  = 1;
  ram[12733]  = 1;
  ram[12734]  = 1;
  ram[12735]  = 1;
  ram[12736]  = 1;
  ram[12737]  = 1;
  ram[12738]  = 1;
  ram[12739]  = 1;
  ram[12740]  = 1;
  ram[12741]  = 1;
  ram[12742]  = 1;
  ram[12743]  = 1;
  ram[12744]  = 1;
  ram[12745]  = 1;
  ram[12746]  = 1;
  ram[12747]  = 1;
  ram[12748]  = 1;
  ram[12749]  = 1;
  ram[12750]  = 1;
  ram[12751]  = 1;
  ram[12752]  = 1;
  ram[12753]  = 1;
  ram[12754]  = 1;
  ram[12755]  = 1;
  ram[12756]  = 1;
  ram[12757]  = 1;
  ram[12758]  = 1;
  ram[12759]  = 1;
  ram[12760]  = 1;
  ram[12761]  = 1;
  ram[12762]  = 1;
  ram[12763]  = 1;
  ram[12764]  = 1;
  ram[12765]  = 1;
  ram[12766]  = 1;
  ram[12767]  = 1;
  ram[12768]  = 1;
  ram[12769]  = 1;
  ram[12770]  = 1;
  ram[12771]  = 1;
  ram[12772]  = 1;
  ram[12773]  = 1;
  ram[12774]  = 1;
  ram[12775]  = 1;
  ram[12776]  = 1;
  ram[12777]  = 1;
  ram[12778]  = 1;
  ram[12779]  = 1;
  ram[12780]  = 1;
  ram[12781]  = 1;
  ram[12782]  = 1;
  ram[12783]  = 1;
  ram[12784]  = 1;
  ram[12785]  = 1;
  ram[12786]  = 1;
  ram[12787]  = 1;
  ram[12788]  = 1;
  ram[12789]  = 1;
  ram[12790]  = 1;
  ram[12791]  = 1;
  ram[12792]  = 1;
  ram[12793]  = 1;
  ram[12794]  = 1;
  ram[12795]  = 1;
  ram[12796]  = 1;
  ram[12797]  = 1;
  ram[12798]  = 1;
  ram[12799]  = 1;
  ram[12800]  = 1;
  ram[12801]  = 1;
  ram[12802]  = 1;
  ram[12803]  = 1;
  ram[12804]  = 1;
  ram[12805]  = 1;
  ram[12806]  = 1;
  ram[12807]  = 1;
  ram[12808]  = 1;
  ram[12809]  = 1;
  ram[12810]  = 1;
  ram[12811]  = 1;
  ram[12812]  = 1;
  ram[12813]  = 1;
  ram[12814]  = 1;
  ram[12815]  = 1;
  ram[12816]  = 1;
  ram[12817]  = 1;
  ram[12818]  = 1;
  ram[12819]  = 1;
  ram[12820]  = 1;
  ram[12821]  = 1;
  ram[12822]  = 1;
  ram[12823]  = 1;
  ram[12824]  = 1;
  ram[12825]  = 1;
  ram[12826]  = 1;
  ram[12827]  = 1;
  ram[12828]  = 1;
  ram[12829]  = 1;
  ram[12830]  = 1;
  ram[12831]  = 1;
  ram[12832]  = 1;
  ram[12833]  = 1;
  ram[12834]  = 1;
  ram[12835]  = 1;
  ram[12836]  = 1;
  ram[12837]  = 1;
  ram[12838]  = 1;
  ram[12839]  = 1;
  ram[12840]  = 1;
  ram[12841]  = 1;
  ram[12842]  = 1;
  ram[12843]  = 1;
  ram[12844]  = 1;
  ram[12845]  = 1;
  ram[12846]  = 1;
  ram[12847]  = 1;
  ram[12848]  = 1;
  ram[12849]  = 1;
  ram[12850]  = 1;
  ram[12851]  = 1;
  ram[12852]  = 1;
  ram[12853]  = 1;
  ram[12854]  = 1;
  ram[12855]  = 1;
  ram[12856]  = 1;
  ram[12857]  = 1;
  ram[12858]  = 1;
  ram[12859]  = 1;
  ram[12860]  = 1;
  ram[12861]  = 1;
  ram[12862]  = 1;
  ram[12863]  = 1;
  ram[12864]  = 1;
  ram[12865]  = 1;
  ram[12866]  = 1;
  ram[12867]  = 1;
  ram[12868]  = 1;
  ram[12869]  = 1;
  ram[12870]  = 1;
  ram[12871]  = 1;
  ram[12872]  = 1;
  ram[12873]  = 1;
  ram[12874]  = 1;
  ram[12875]  = 1;
  ram[12876]  = 1;
  ram[12877]  = 1;
  ram[12878]  = 1;
  ram[12879]  = 1;
  ram[12880]  = 1;
  ram[12881]  = 1;
  ram[12882]  = 1;
  ram[12883]  = 1;
  ram[12884]  = 1;
  ram[12885]  = 1;
  ram[12886]  = 1;
  ram[12887]  = 1;
  ram[12888]  = 1;
  ram[12889]  = 1;
  ram[12890]  = 1;
  ram[12891]  = 1;
  ram[12892]  = 1;
  ram[12893]  = 1;
  ram[12894]  = 1;
  ram[12895]  = 1;
  ram[12896]  = 1;
  ram[12897]  = 1;
  ram[12898]  = 1;
  ram[12899]  = 1;
  ram[12900]  = 1;
  ram[12901]  = 1;
  ram[12902]  = 1;
  ram[12903]  = 1;
  ram[12904]  = 1;
  ram[12905]  = 1;
  ram[12906]  = 1;
  ram[12907]  = 1;
  ram[12908]  = 1;
  ram[12909]  = 1;
  ram[12910]  = 1;
  ram[12911]  = 1;
  ram[12912]  = 1;
  ram[12913]  = 1;
  ram[12914]  = 1;
  ram[12915]  = 1;
  ram[12916]  = 1;
  ram[12917]  = 1;
  ram[12918]  = 1;
  ram[12919]  = 1;
  ram[12920]  = 1;
  ram[12921]  = 1;
  ram[12922]  = 1;
  ram[12923]  = 1;
  ram[12924]  = 1;
  ram[12925]  = 1;
  ram[12926]  = 1;
  ram[12927]  = 1;
  ram[12928]  = 1;
  ram[12929]  = 1;
  ram[12930]  = 1;
  ram[12931]  = 1;
  ram[12932]  = 1;
  ram[12933]  = 1;
  ram[12934]  = 1;
  ram[12935]  = 1;
  ram[12936]  = 1;
  ram[12937]  = 1;
  ram[12938]  = 1;
  ram[12939]  = 1;
  ram[12940]  = 1;
  ram[12941]  = 1;
  ram[12942]  = 1;
  ram[12943]  = 1;
  ram[12944]  = 1;
  ram[12945]  = 1;
  ram[12946]  = 1;
  ram[12947]  = 1;
  ram[12948]  = 1;
  ram[12949]  = 1;
  ram[12950]  = 1;
  ram[12951]  = 1;
  ram[12952]  = 1;
  ram[12953]  = 1;
  ram[12954]  = 1;
  ram[12955]  = 1;
  ram[12956]  = 1;
  ram[12957]  = 1;
  ram[12958]  = 1;
  ram[12959]  = 1;
  ram[12960]  = 1;
  ram[12961]  = 1;
  ram[12962]  = 1;
  ram[12963]  = 1;
  ram[12964]  = 1;
  ram[12965]  = 1;
  ram[12966]  = 1;
  ram[12967]  = 1;
  ram[12968]  = 1;
  ram[12969]  = 1;
  ram[12970]  = 1;
  ram[12971]  = 1;
  ram[12972]  = 1;
  ram[12973]  = 1;
  ram[12974]  = 1;
  ram[12975]  = 1;
  ram[12976]  = 1;
  ram[12977]  = 1;
  ram[12978]  = 1;
  ram[12979]  = 1;
  ram[12980]  = 1;
  ram[12981]  = 1;
  ram[12982]  = 1;
  ram[12983]  = 1;
  ram[12984]  = 1;
  ram[12985]  = 1;
  ram[12986]  = 1;
  ram[12987]  = 1;
  ram[12988]  = 1;
  ram[12989]  = 1;
  ram[12990]  = 1;
  ram[12991]  = 1;
  ram[12992]  = 1;
  ram[12993]  = 1;
  ram[12994]  = 1;
  ram[12995]  = 1;
  ram[12996]  = 1;
  ram[12997]  = 1;
  ram[12998]  = 1;
  ram[12999]  = 1;
  ram[13000]  = 1;
  ram[13001]  = 1;
  ram[13002]  = 1;
  ram[13003]  = 1;
  ram[13004]  = 1;
  ram[13005]  = 1;
  ram[13006]  = 1;
  ram[13007]  = 1;
  ram[13008]  = 1;
  ram[13009]  = 1;
  ram[13010]  = 1;
  ram[13011]  = 1;
  ram[13012]  = 1;
  ram[13013]  = 1;
  ram[13014]  = 1;
  ram[13015]  = 1;
  ram[13016]  = 1;
  ram[13017]  = 1;
  ram[13018]  = 1;
  ram[13019]  = 1;
  ram[13020]  = 1;
  ram[13021]  = 1;
  ram[13022]  = 1;
  ram[13023]  = 1;
  ram[13024]  = 1;
  ram[13025]  = 1;
  ram[13026]  = 1;
  ram[13027]  = 1;
  ram[13028]  = 1;
  ram[13029]  = 1;
  ram[13030]  = 1;
  ram[13031]  = 1;
  ram[13032]  = 1;
  ram[13033]  = 1;
  ram[13034]  = 1;
  ram[13035]  = 1;
  ram[13036]  = 1;
  ram[13037]  = 1;
  ram[13038]  = 1;
  ram[13039]  = 1;
  ram[13040]  = 1;
  ram[13041]  = 1;
  ram[13042]  = 1;
  ram[13043]  = 1;
  ram[13044]  = 1;
  ram[13045]  = 1;
  ram[13046]  = 1;
  ram[13047]  = 1;
  ram[13048]  = 1;
  ram[13049]  = 1;
  ram[13050]  = 1;
  ram[13051]  = 1;
  ram[13052]  = 1;
  ram[13053]  = 1;
  ram[13054]  = 1;
  ram[13055]  = 1;
  ram[13056]  = 1;
  ram[13057]  = 1;
  ram[13058]  = 1;
  ram[13059]  = 1;
  ram[13060]  = 1;
  ram[13061]  = 1;
  ram[13062]  = 1;
  ram[13063]  = 1;
  ram[13064]  = 1;
  ram[13065]  = 1;
  ram[13066]  = 1;
  ram[13067]  = 1;
  ram[13068]  = 1;
  ram[13069]  = 1;
  ram[13070]  = 1;
  ram[13071]  = 1;
  ram[13072]  = 1;
  ram[13073]  = 1;
  ram[13074]  = 1;
  ram[13075]  = 1;
  ram[13076]  = 1;
  ram[13077]  = 1;
  ram[13078]  = 1;
  ram[13079]  = 1;
  ram[13080]  = 1;
  ram[13081]  = 1;
  ram[13082]  = 1;
  ram[13083]  = 1;
  ram[13084]  = 1;
  ram[13085]  = 1;
  ram[13086]  = 1;
  ram[13087]  = 1;
  ram[13088]  = 1;
  ram[13089]  = 1;
  ram[13090]  = 1;
  ram[13091]  = 1;
  ram[13092]  = 1;
  ram[13093]  = 1;
  ram[13094]  = 1;
  ram[13095]  = 1;
  ram[13096]  = 1;
  ram[13097]  = 1;
  ram[13098]  = 1;
  ram[13099]  = 1;
  ram[13100]  = 1;
  ram[13101]  = 1;
  ram[13102]  = 1;
  ram[13103]  = 1;
  ram[13104]  = 1;
  ram[13105]  = 1;
  ram[13106]  = 1;
  ram[13107]  = 1;
  ram[13108]  = 1;
  ram[13109]  = 1;
  ram[13110]  = 1;
  ram[13111]  = 1;
  ram[13112]  = 1;
  ram[13113]  = 1;
  ram[13114]  = 1;
  ram[13115]  = 1;
  ram[13116]  = 1;
  ram[13117]  = 1;
  ram[13118]  = 1;
  ram[13119]  = 1;
  ram[13120]  = 1;
  ram[13121]  = 1;
  ram[13122]  = 1;
  ram[13123]  = 1;
  ram[13124]  = 1;
  ram[13125]  = 1;
  ram[13126]  = 1;
  ram[13127]  = 1;
  ram[13128]  = 1;
  ram[13129]  = 1;
  ram[13130]  = 1;
  ram[13131]  = 1;
  ram[13132]  = 1;
  ram[13133]  = 1;
  ram[13134]  = 1;
  ram[13135]  = 1;
  ram[13136]  = 1;
  ram[13137]  = 1;
  ram[13138]  = 1;
  ram[13139]  = 1;
  ram[13140]  = 1;
  ram[13141]  = 1;
  ram[13142]  = 1;
  ram[13143]  = 1;
  ram[13144]  = 1;
  ram[13145]  = 1;
  ram[13146]  = 1;
  ram[13147]  = 1;
  ram[13148]  = 1;
  ram[13149]  = 1;
  ram[13150]  = 1;
  ram[13151]  = 1;
  ram[13152]  = 1;
  ram[13153]  = 1;
  ram[13154]  = 1;
  ram[13155]  = 1;
  ram[13156]  = 1;
  ram[13157]  = 1;
  ram[13158]  = 1;
  ram[13159]  = 1;
  ram[13160]  = 1;
  ram[13161]  = 1;
  ram[13162]  = 1;
  ram[13163]  = 1;
  ram[13164]  = 1;
  ram[13165]  = 1;
  ram[13166]  = 1;
  ram[13167]  = 1;
  ram[13168]  = 1;
  ram[13169]  = 1;
  ram[13170]  = 1;
  ram[13171]  = 1;
  ram[13172]  = 1;
  ram[13173]  = 1;
  ram[13174]  = 1;
  ram[13175]  = 1;
  ram[13176]  = 1;
  ram[13177]  = 1;
  ram[13178]  = 1;
  ram[13179]  = 1;
  ram[13180]  = 1;
  ram[13181]  = 1;
  ram[13182]  = 1;
  ram[13183]  = 1;
  ram[13184]  = 1;
  ram[13185]  = 1;
  ram[13186]  = 1;
  ram[13187]  = 1;
  ram[13188]  = 1;
  ram[13189]  = 1;
  ram[13190]  = 1;
  ram[13191]  = 1;
  ram[13192]  = 1;
  ram[13193]  = 1;
  ram[13194]  = 1;
  ram[13195]  = 1;
  ram[13196]  = 1;
  ram[13197]  = 1;
  ram[13198]  = 1;
  ram[13199]  = 1;
  ram[13200]  = 1;
  ram[13201]  = 1;
  ram[13202]  = 1;
  ram[13203]  = 1;
  ram[13204]  = 1;
  ram[13205]  = 1;
  ram[13206]  = 1;
  ram[13207]  = 1;
  ram[13208]  = 1;
  ram[13209]  = 1;
  ram[13210]  = 1;
  ram[13211]  = 1;
  ram[13212]  = 1;
  ram[13213]  = 1;
  ram[13214]  = 1;
  ram[13215]  = 1;
  ram[13216]  = 1;
  ram[13217]  = 1;
  ram[13218]  = 1;
  ram[13219]  = 1;
  ram[13220]  = 1;
  ram[13221]  = 1;
  ram[13222]  = 1;
  ram[13223]  = 1;
  ram[13224]  = 1;
  ram[13225]  = 1;
  ram[13226]  = 1;
  ram[13227]  = 1;
  ram[13228]  = 1;
  ram[13229]  = 1;
  ram[13230]  = 1;
  ram[13231]  = 1;
  ram[13232]  = 1;
  ram[13233]  = 1;
  ram[13234]  = 1;
  ram[13235]  = 1;
  ram[13236]  = 1;
  ram[13237]  = 1;
  ram[13238]  = 1;
  ram[13239]  = 1;
  ram[13240]  = 1;
  ram[13241]  = 1;
  ram[13242]  = 1;
  ram[13243]  = 1;
  ram[13244]  = 1;
  ram[13245]  = 1;
  ram[13246]  = 1;
  ram[13247]  = 1;
  ram[13248]  = 1;
  ram[13249]  = 1;
  ram[13250]  = 1;
  ram[13251]  = 1;
  ram[13252]  = 1;
  ram[13253]  = 1;
  ram[13254]  = 1;
  ram[13255]  = 1;
  ram[13256]  = 1;
  ram[13257]  = 1;
  ram[13258]  = 1;
  ram[13259]  = 1;
  ram[13260]  = 1;
  ram[13261]  = 1;
  ram[13262]  = 1;
  ram[13263]  = 1;
  ram[13264]  = 1;
  ram[13265]  = 1;
  ram[13266]  = 1;
  ram[13267]  = 1;
  ram[13268]  = 1;
  ram[13269]  = 1;
  ram[13270]  = 1;
  ram[13271]  = 1;
  ram[13272]  = 1;
  ram[13273]  = 1;
  ram[13274]  = 1;
  ram[13275]  = 1;
  ram[13276]  = 1;
  ram[13277]  = 1;
  ram[13278]  = 1;
  ram[13279]  = 1;
  ram[13280]  = 1;
  ram[13281]  = 1;
  ram[13282]  = 1;
  ram[13283]  = 1;
  ram[13284]  = 1;
  ram[13285]  = 1;
  ram[13286]  = 1;
  ram[13287]  = 1;
  ram[13288]  = 1;
  ram[13289]  = 1;
  ram[13290]  = 1;
  ram[13291]  = 1;
  ram[13292]  = 1;
  ram[13293]  = 1;
  ram[13294]  = 1;
  ram[13295]  = 1;
  ram[13296]  = 1;
  ram[13297]  = 1;
  ram[13298]  = 1;
  ram[13299]  = 1;
  ram[13300]  = 1;
  ram[13301]  = 1;
  ram[13302]  = 1;
  ram[13303]  = 1;
  ram[13304]  = 1;
  ram[13305]  = 1;
  ram[13306]  = 1;
  ram[13307]  = 1;
  ram[13308]  = 1;
  ram[13309]  = 1;
  ram[13310]  = 1;
  ram[13311]  = 1;
  ram[13312]  = 1;
  ram[13313]  = 1;
  ram[13314]  = 1;
  ram[13315]  = 1;
  ram[13316]  = 1;
  ram[13317]  = 1;
  ram[13318]  = 1;
  ram[13319]  = 1;
  ram[13320]  = 1;
  ram[13321]  = 1;
  ram[13322]  = 1;
  ram[13323]  = 1;
  ram[13324]  = 1;
  ram[13325]  = 1;
  ram[13326]  = 1;
  ram[13327]  = 1;
  ram[13328]  = 1;
  ram[13329]  = 1;
  ram[13330]  = 1;
  ram[13331]  = 1;
  ram[13332]  = 1;
  ram[13333]  = 1;
  ram[13334]  = 1;
  ram[13335]  = 1;
  ram[13336]  = 1;
  ram[13337]  = 1;
  ram[13338]  = 1;
  ram[13339]  = 1;
  ram[13340]  = 1;
  ram[13341]  = 1;
  ram[13342]  = 1;
  ram[13343]  = 1;
  ram[13344]  = 1;
  ram[13345]  = 1;
  ram[13346]  = 1;
  ram[13347]  = 1;
  ram[13348]  = 1;
  ram[13349]  = 1;
  ram[13350]  = 1;
  ram[13351]  = 1;
  ram[13352]  = 1;
  ram[13353]  = 1;
  ram[13354]  = 1;
  ram[13355]  = 1;
  ram[13356]  = 1;
  ram[13357]  = 1;
  ram[13358]  = 1;
  ram[13359]  = 1;
  ram[13360]  = 1;
  ram[13361]  = 1;
  ram[13362]  = 1;
  ram[13363]  = 1;
  ram[13364]  = 1;
  ram[13365]  = 1;
  ram[13366]  = 1;
  ram[13367]  = 1;
  ram[13368]  = 1;
  ram[13369]  = 1;
  ram[13370]  = 1;
  ram[13371]  = 1;
  ram[13372]  = 1;
  ram[13373]  = 1;
  ram[13374]  = 1;
  ram[13375]  = 1;
  ram[13376]  = 1;
  ram[13377]  = 1;
  ram[13378]  = 1;
  ram[13379]  = 1;
  ram[13380]  = 1;
  ram[13381]  = 1;
  ram[13382]  = 1;
  ram[13383]  = 1;
  ram[13384]  = 1;
  ram[13385]  = 1;
  ram[13386]  = 1;
  ram[13387]  = 1;
  ram[13388]  = 1;
  ram[13389]  = 1;
  ram[13390]  = 1;
  ram[13391]  = 1;
  ram[13392]  = 1;
  ram[13393]  = 1;
  ram[13394]  = 1;
  ram[13395]  = 1;
  ram[13396]  = 1;
  ram[13397]  = 1;
  ram[13398]  = 1;
  ram[13399]  = 1;
  ram[13400]  = 1;
  ram[13401]  = 1;
  ram[13402]  = 1;
  ram[13403]  = 1;
  ram[13404]  = 1;
  ram[13405]  = 1;
  ram[13406]  = 1;
  ram[13407]  = 1;
  ram[13408]  = 1;
  ram[13409]  = 1;
  ram[13410]  = 1;
  ram[13411]  = 1;
  ram[13412]  = 1;
  ram[13413]  = 1;
  ram[13414]  = 1;
  ram[13415]  = 1;
  ram[13416]  = 1;
  ram[13417]  = 1;
  ram[13418]  = 1;
  ram[13419]  = 1;
  ram[13420]  = 1;
  ram[13421]  = 1;
  ram[13422]  = 1;
  ram[13423]  = 1;
  ram[13424]  = 1;
  ram[13425]  = 1;
  ram[13426]  = 1;
  ram[13427]  = 1;
  ram[13428]  = 1;
  ram[13429]  = 1;
  ram[13430]  = 1;
  ram[13431]  = 1;
  ram[13432]  = 1;
  ram[13433]  = 1;
  ram[13434]  = 1;
  ram[13435]  = 1;
  ram[13436]  = 1;
  ram[13437]  = 1;
  ram[13438]  = 1;
  ram[13439]  = 1;
  ram[13440]  = 1;
  ram[13441]  = 1;
  ram[13442]  = 1;
  ram[13443]  = 1;
  ram[13444]  = 1;
  ram[13445]  = 1;
  ram[13446]  = 1;
  ram[13447]  = 1;
  ram[13448]  = 1;
  ram[13449]  = 1;
  ram[13450]  = 1;
  ram[13451]  = 1;
  ram[13452]  = 1;
  ram[13453]  = 1;
  ram[13454]  = 1;
  ram[13455]  = 1;
  ram[13456]  = 1;
  ram[13457]  = 1;
  ram[13458]  = 1;
  ram[13459]  = 1;
  ram[13460]  = 1;
  ram[13461]  = 1;
  ram[13462]  = 1;
  ram[13463]  = 1;
  ram[13464]  = 1;
  ram[13465]  = 1;
  ram[13466]  = 1;
  ram[13467]  = 1;
  ram[13468]  = 1;
  ram[13469]  = 1;
  ram[13470]  = 1;
  ram[13471]  = 1;
  ram[13472]  = 1;
  ram[13473]  = 1;
  ram[13474]  = 1;
  ram[13475]  = 1;
  ram[13476]  = 1;
  ram[13477]  = 1;
  ram[13478]  = 1;
  ram[13479]  = 1;
  ram[13480]  = 1;
  ram[13481]  = 1;
  ram[13482]  = 1;
  ram[13483]  = 1;
  ram[13484]  = 1;
  ram[13485]  = 1;
  ram[13486]  = 1;
  ram[13487]  = 1;
  ram[13488]  = 1;
  ram[13489]  = 1;
  ram[13490]  = 1;
  ram[13491]  = 1;
  ram[13492]  = 1;
  ram[13493]  = 1;
  ram[13494]  = 1;
  ram[13495]  = 1;
  ram[13496]  = 1;
  ram[13497]  = 1;
  ram[13498]  = 1;
  ram[13499]  = 1;
  ram[13500]  = 1;
  ram[13501]  = 1;
  ram[13502]  = 1;
  ram[13503]  = 1;
  ram[13504]  = 1;
  ram[13505]  = 1;
  ram[13506]  = 1;
  ram[13507]  = 1;
  ram[13508]  = 1;
  ram[13509]  = 1;
  ram[13510]  = 1;
  ram[13511]  = 1;
  ram[13512]  = 1;
  ram[13513]  = 1;
  ram[13514]  = 1;
  ram[13515]  = 1;
  ram[13516]  = 1;
  ram[13517]  = 1;
  ram[13518]  = 1;
  ram[13519]  = 1;
  ram[13520]  = 1;
  ram[13521]  = 1;
  ram[13522]  = 1;
  ram[13523]  = 1;
  ram[13524]  = 1;
  ram[13525]  = 1;
  ram[13526]  = 1;
  ram[13527]  = 1;
  ram[13528]  = 1;
  ram[13529]  = 1;
  ram[13530]  = 1;
  ram[13531]  = 1;
  ram[13532]  = 1;
  ram[13533]  = 1;
  ram[13534]  = 1;
  ram[13535]  = 1;
  ram[13536]  = 1;
  ram[13537]  = 1;
  ram[13538]  = 1;
  ram[13539]  = 1;
  ram[13540]  = 1;
  ram[13541]  = 1;
  ram[13542]  = 1;
  ram[13543]  = 1;
  ram[13544]  = 1;
  ram[13545]  = 1;
  ram[13546]  = 1;
  ram[13547]  = 1;
  ram[13548]  = 1;
  ram[13549]  = 1;
  ram[13550]  = 1;
  ram[13551]  = 1;
  ram[13552]  = 1;
  ram[13553]  = 1;
  ram[13554]  = 1;
  ram[13555]  = 1;
  ram[13556]  = 1;
  ram[13557]  = 1;
  ram[13558]  = 1;
  ram[13559]  = 1;
  ram[13560]  = 1;
  ram[13561]  = 1;
  ram[13562]  = 1;
  ram[13563]  = 1;
  ram[13564]  = 1;
  ram[13565]  = 1;
  ram[13566]  = 1;
  ram[13567]  = 1;
  ram[13568]  = 1;
  ram[13569]  = 1;
  ram[13570]  = 1;
  ram[13571]  = 1;
  ram[13572]  = 1;
  ram[13573]  = 1;
  ram[13574]  = 1;
  ram[13575]  = 1;
  ram[13576]  = 1;
  ram[13577]  = 1;
  ram[13578]  = 1;
  ram[13579]  = 1;
  ram[13580]  = 1;
  ram[13581]  = 1;
  ram[13582]  = 1;
  ram[13583]  = 1;
  ram[13584]  = 1;
  ram[13585]  = 1;
  ram[13586]  = 1;
  ram[13587]  = 1;
  ram[13588]  = 1;
  ram[13589]  = 1;
  ram[13590]  = 1;
  ram[13591]  = 1;
  ram[13592]  = 1;
  ram[13593]  = 1;
  ram[13594]  = 1;
  ram[13595]  = 1;
  ram[13596]  = 1;
  ram[13597]  = 1;
  ram[13598]  = 1;
  ram[13599]  = 1;
  ram[13600]  = 1;
  ram[13601]  = 1;
  ram[13602]  = 1;
  ram[13603]  = 1;
  ram[13604]  = 1;
  ram[13605]  = 1;
  ram[13606]  = 1;
  ram[13607]  = 1;
  ram[13608]  = 1;
  ram[13609]  = 1;
  ram[13610]  = 1;
  ram[13611]  = 1;
  ram[13612]  = 1;
  ram[13613]  = 1;
  ram[13614]  = 1;
  ram[13615]  = 1;
  ram[13616]  = 1;
  ram[13617]  = 1;
  ram[13618]  = 1;
  ram[13619]  = 1;
  ram[13620]  = 1;
  ram[13621]  = 1;
  ram[13622]  = 1;
  ram[13623]  = 1;
  ram[13624]  = 1;
  ram[13625]  = 1;
  ram[13626]  = 1;
  ram[13627]  = 1;
  ram[13628]  = 1;
  ram[13629]  = 1;
  ram[13630]  = 1;
  ram[13631]  = 1;
  ram[13632]  = 1;
  ram[13633]  = 1;
  ram[13634]  = 1;
  ram[13635]  = 1;
  ram[13636]  = 1;
  ram[13637]  = 1;
  ram[13638]  = 1;
  ram[13639]  = 1;
  ram[13640]  = 1;
  ram[13641]  = 1;
  ram[13642]  = 1;
  ram[13643]  = 1;
  ram[13644]  = 1;
  ram[13645]  = 1;
  ram[13646]  = 1;
  ram[13647]  = 1;
  ram[13648]  = 1;
  ram[13649]  = 1;
  ram[13650]  = 1;
  ram[13651]  = 1;
  ram[13652]  = 1;
  ram[13653]  = 1;
  ram[13654]  = 1;
  ram[13655]  = 1;
  ram[13656]  = 1;
  ram[13657]  = 1;
  ram[13658]  = 1;
  ram[13659]  = 1;
  ram[13660]  = 1;
  ram[13661]  = 1;
  ram[13662]  = 1;
  ram[13663]  = 1;
  ram[13664]  = 1;
  ram[13665]  = 1;
  ram[13666]  = 1;
  ram[13667]  = 1;
  ram[13668]  = 1;
  ram[13669]  = 1;
  ram[13670]  = 1;
  ram[13671]  = 1;
  ram[13672]  = 1;
  ram[13673]  = 1;
  ram[13674]  = 1;
  ram[13675]  = 1;
  ram[13676]  = 1;
  ram[13677]  = 1;
  ram[13678]  = 1;
  ram[13679]  = 1;
  ram[13680]  = 1;
  ram[13681]  = 1;
  ram[13682]  = 1;
  ram[13683]  = 1;
  ram[13684]  = 1;
  ram[13685]  = 1;
  ram[13686]  = 1;
  ram[13687]  = 1;
  ram[13688]  = 1;
  ram[13689]  = 1;
  ram[13690]  = 1;
  ram[13691]  = 1;
  ram[13692]  = 1;
  ram[13693]  = 1;
  ram[13694]  = 1;
  ram[13695]  = 1;
  ram[13696]  = 1;
  ram[13697]  = 1;
  ram[13698]  = 1;
  ram[13699]  = 1;
  ram[13700]  = 1;
  ram[13701]  = 1;
  ram[13702]  = 1;
  ram[13703]  = 1;
  ram[13704]  = 1;
  ram[13705]  = 1;
  ram[13706]  = 1;
  ram[13707]  = 1;
  ram[13708]  = 1;
  ram[13709]  = 1;
  ram[13710]  = 1;
  ram[13711]  = 1;
  ram[13712]  = 1;
  ram[13713]  = 1;
  ram[13714]  = 1;
  ram[13715]  = 1;
  ram[13716]  = 1;
  ram[13717]  = 1;
  ram[13718]  = 1;
  ram[13719]  = 1;
  ram[13720]  = 1;
  ram[13721]  = 1;
  ram[13722]  = 1;
  ram[13723]  = 1;
  ram[13724]  = 1;
  ram[13725]  = 1;
  ram[13726]  = 1;
  ram[13727]  = 1;
  ram[13728]  = 1;
  ram[13729]  = 1;
  ram[13730]  = 1;
  ram[13731]  = 1;
  ram[13732]  = 1;
  ram[13733]  = 1;
  ram[13734]  = 1;
  ram[13735]  = 1;
  ram[13736]  = 1;
  ram[13737]  = 1;
  ram[13738]  = 1;
  ram[13739]  = 1;
  ram[13740]  = 1;
  ram[13741]  = 1;
  ram[13742]  = 1;
  ram[13743]  = 1;
  ram[13744]  = 1;
  ram[13745]  = 1;
  ram[13746]  = 1;
  ram[13747]  = 1;
  ram[13748]  = 1;
  ram[13749]  = 1;
  ram[13750]  = 1;
  ram[13751]  = 1;
  ram[13752]  = 1;
  ram[13753]  = 1;
  ram[13754]  = 1;
  ram[13755]  = 1;
  ram[13756]  = 1;
  ram[13757]  = 1;
  ram[13758]  = 1;
  ram[13759]  = 1;
  ram[13760]  = 1;
  ram[13761]  = 1;
  ram[13762]  = 1;
  ram[13763]  = 1;
  ram[13764]  = 1;
  ram[13765]  = 1;
  ram[13766]  = 1;
  ram[13767]  = 1;
  ram[13768]  = 1;
  ram[13769]  = 1;
  ram[13770]  = 1;
  ram[13771]  = 1;
  ram[13772]  = 1;
  ram[13773]  = 1;
  ram[13774]  = 1;
  ram[13775]  = 1;
  ram[13776]  = 1;
  ram[13777]  = 1;
  ram[13778]  = 1;
  ram[13779]  = 1;
  ram[13780]  = 1;
  ram[13781]  = 1;
  ram[13782]  = 1;
  ram[13783]  = 1;
  ram[13784]  = 1;
  ram[13785]  = 1;
  ram[13786]  = 1;
  ram[13787]  = 1;
  ram[13788]  = 1;
  ram[13789]  = 1;
  ram[13790]  = 1;
  ram[13791]  = 1;
  ram[13792]  = 1;
  ram[13793]  = 1;
  ram[13794]  = 1;
  ram[13795]  = 1;
  ram[13796]  = 1;
  ram[13797]  = 1;
  ram[13798]  = 1;
  ram[13799]  = 1;
  ram[13800]  = 1;
  ram[13801]  = 1;
  ram[13802]  = 1;
  ram[13803]  = 1;
  ram[13804]  = 1;
  ram[13805]  = 1;
  ram[13806]  = 1;
  ram[13807]  = 1;
  ram[13808]  = 1;
  ram[13809]  = 1;
  ram[13810]  = 1;
  ram[13811]  = 1;
  ram[13812]  = 1;
  ram[13813]  = 1;
  ram[13814]  = 1;
  ram[13815]  = 1;
  ram[13816]  = 1;
  ram[13817]  = 1;
  ram[13818]  = 1;
  ram[13819]  = 1;
  ram[13820]  = 1;
  ram[13821]  = 1;
  ram[13822]  = 1;
  ram[13823]  = 1;
  ram[13824]  = 1;
  ram[13825]  = 1;
  ram[13826]  = 1;
  ram[13827]  = 1;
  ram[13828]  = 1;
  ram[13829]  = 1;
  ram[13830]  = 1;
  ram[13831]  = 1;
  ram[13832]  = 1;
  ram[13833]  = 1;
  ram[13834]  = 1;
  ram[13835]  = 1;
  ram[13836]  = 1;
  ram[13837]  = 1;
  ram[13838]  = 1;
  ram[13839]  = 1;
  ram[13840]  = 1;
  ram[13841]  = 1;
  ram[13842]  = 1;
  ram[13843]  = 1;
  ram[13844]  = 1;
  ram[13845]  = 1;
  ram[13846]  = 1;
  ram[13847]  = 1;
  ram[13848]  = 1;
  ram[13849]  = 1;
  ram[13850]  = 1;
  ram[13851]  = 1;
  ram[13852]  = 1;
  ram[13853]  = 1;
  ram[13854]  = 1;
  ram[13855]  = 1;
  ram[13856]  = 1;
  ram[13857]  = 1;
  ram[13858]  = 1;
  ram[13859]  = 1;
  ram[13860]  = 1;
  ram[13861]  = 1;
  ram[13862]  = 1;
  ram[13863]  = 1;
  ram[13864]  = 1;
  ram[13865]  = 1;
  ram[13866]  = 1;
  ram[13867]  = 1;
  ram[13868]  = 1;
  ram[13869]  = 1;
  ram[13870]  = 1;
  ram[13871]  = 1;
  ram[13872]  = 1;
  ram[13873]  = 1;
  ram[13874]  = 1;
  ram[13875]  = 1;
  ram[13876]  = 1;
  ram[13877]  = 1;
  ram[13878]  = 1;
  ram[13879]  = 1;
  ram[13880]  = 1;
  ram[13881]  = 1;
  ram[13882]  = 1;
  ram[13883]  = 1;
  ram[13884]  = 1;
  ram[13885]  = 1;
  ram[13886]  = 1;
  ram[13887]  = 1;
  ram[13888]  = 1;
  ram[13889]  = 1;
  ram[13890]  = 1;
  ram[13891]  = 1;
  ram[13892]  = 1;
  ram[13893]  = 1;
  ram[13894]  = 1;
  ram[13895]  = 1;
  ram[13896]  = 1;
  ram[13897]  = 1;
  ram[13898]  = 1;
  ram[13899]  = 1;
  ram[13900]  = 1;
  ram[13901]  = 1;
  ram[13902]  = 1;
  ram[13903]  = 1;
  ram[13904]  = 1;
  ram[13905]  = 1;
  ram[13906]  = 1;
  ram[13907]  = 1;
  ram[13908]  = 1;
  ram[13909]  = 1;
  ram[13910]  = 1;
  ram[13911]  = 1;
  ram[13912]  = 1;
  ram[13913]  = 1;
  ram[13914]  = 1;
  ram[13915]  = 1;
  ram[13916]  = 1;
  ram[13917]  = 1;
  ram[13918]  = 1;
  ram[13919]  = 1;
  ram[13920]  = 1;
  ram[13921]  = 1;
  ram[13922]  = 1;
  ram[13923]  = 1;
  ram[13924]  = 1;
  ram[13925]  = 1;
  ram[13926]  = 1;
  ram[13927]  = 1;
  ram[13928]  = 1;
  ram[13929]  = 1;
  ram[13930]  = 1;
  ram[13931]  = 1;
  ram[13932]  = 1;
  ram[13933]  = 1;
  ram[13934]  = 1;
  ram[13935]  = 1;
  ram[13936]  = 1;
  ram[13937]  = 1;
  ram[13938]  = 1;
  ram[13939]  = 1;
  ram[13940]  = 1;
  ram[13941]  = 1;
  ram[13942]  = 1;
  ram[13943]  = 1;
  ram[13944]  = 1;
  ram[13945]  = 1;
  ram[13946]  = 1;
  ram[13947]  = 1;
  ram[13948]  = 1;
  ram[13949]  = 1;
  ram[13950]  = 1;
  ram[13951]  = 1;
  ram[13952]  = 1;
  ram[13953]  = 1;
  ram[13954]  = 1;
  ram[13955]  = 1;
  ram[13956]  = 1;
  ram[13957]  = 1;
  ram[13958]  = 1;
  ram[13959]  = 1;
  ram[13960]  = 1;
  ram[13961]  = 1;
  ram[13962]  = 1;
  ram[13963]  = 1;
  ram[13964]  = 1;
  ram[13965]  = 1;
  ram[13966]  = 1;
  ram[13967]  = 1;
  ram[13968]  = 1;
  ram[13969]  = 1;
  ram[13970]  = 1;
  ram[13971]  = 1;
  ram[13972]  = 1;
  ram[13973]  = 1;
  ram[13974]  = 1;
  ram[13975]  = 1;
  ram[13976]  = 1;
  ram[13977]  = 1;
  ram[13978]  = 1;
  ram[13979]  = 1;
  ram[13980]  = 1;
  ram[13981]  = 1;
  ram[13982]  = 1;
  ram[13983]  = 1;
  ram[13984]  = 1;
  ram[13985]  = 1;
  ram[13986]  = 1;
  ram[13987]  = 1;
  ram[13988]  = 1;
  ram[13989]  = 1;
  ram[13990]  = 1;
  ram[13991]  = 1;
  ram[13992]  = 1;
  ram[13993]  = 1;
  ram[13994]  = 1;
  ram[13995]  = 1;
  ram[13996]  = 1;
  ram[13997]  = 1;
  ram[13998]  = 1;
  ram[13999]  = 1;
  ram[14000]  = 1;
  ram[14001]  = 1;
  ram[14002]  = 1;
  ram[14003]  = 1;
  ram[14004]  = 1;
  ram[14005]  = 1;
  ram[14006]  = 1;
  ram[14007]  = 1;
  ram[14008]  = 1;
  ram[14009]  = 1;
  ram[14010]  = 1;
  ram[14011]  = 1;
  ram[14012]  = 1;
  ram[14013]  = 1;
  ram[14014]  = 1;
  ram[14015]  = 1;
  ram[14016]  = 1;
  ram[14017]  = 1;
  ram[14018]  = 1;
  ram[14019]  = 1;
  ram[14020]  = 1;
  ram[14021]  = 1;
  ram[14022]  = 1;
  ram[14023]  = 1;
  ram[14024]  = 1;
  ram[14025]  = 1;
  ram[14026]  = 1;
  ram[14027]  = 1;
  ram[14028]  = 1;
  ram[14029]  = 1;
  ram[14030]  = 1;
  ram[14031]  = 1;
  ram[14032]  = 1;
  ram[14033]  = 1;
  ram[14034]  = 1;
  ram[14035]  = 1;
  ram[14036]  = 1;
  ram[14037]  = 1;
  ram[14038]  = 1;
  ram[14039]  = 1;
  ram[14040]  = 1;
  ram[14041]  = 1;
  ram[14042]  = 1;
  ram[14043]  = 1;
  ram[14044]  = 1;
  ram[14045]  = 1;
  ram[14046]  = 1;
  ram[14047]  = 1;
  ram[14048]  = 1;
  ram[14049]  = 1;
  ram[14050]  = 1;
  ram[14051]  = 1;
  ram[14052]  = 1;
  ram[14053]  = 1;
  ram[14054]  = 1;
  ram[14055]  = 1;
  ram[14056]  = 1;
  ram[14057]  = 1;
  ram[14058]  = 1;
  ram[14059]  = 1;
  ram[14060]  = 1;
  ram[14061]  = 1;
  ram[14062]  = 1;
  ram[14063]  = 1;
  ram[14064]  = 1;
  ram[14065]  = 1;
  ram[14066]  = 1;
  ram[14067]  = 1;
  ram[14068]  = 1;
  ram[14069]  = 1;
  ram[14070]  = 1;
  ram[14071]  = 1;
  ram[14072]  = 1;
  ram[14073]  = 1;
  ram[14074]  = 1;
  ram[14075]  = 1;
  ram[14076]  = 1;
  ram[14077]  = 1;
  ram[14078]  = 1;
  ram[14079]  = 1;
  ram[14080]  = 1;
  ram[14081]  = 1;
  ram[14082]  = 1;
  ram[14083]  = 1;
  ram[14084]  = 1;
  ram[14085]  = 1;
  ram[14086]  = 1;
  ram[14087]  = 1;
  ram[14088]  = 1;
  ram[14089]  = 1;
  ram[14090]  = 1;
  ram[14091]  = 1;
  ram[14092]  = 1;
  ram[14093]  = 1;
  ram[14094]  = 1;
  ram[14095]  = 1;
  ram[14096]  = 1;
  ram[14097]  = 1;
  ram[14098]  = 1;
  ram[14099]  = 1;
  ram[14100]  = 1;
  ram[14101]  = 1;
  ram[14102]  = 1;
  ram[14103]  = 1;
  ram[14104]  = 1;
  ram[14105]  = 1;
  ram[14106]  = 1;
  ram[14107]  = 1;
  ram[14108]  = 1;
  ram[14109]  = 1;
  ram[14110]  = 1;
  ram[14111]  = 1;
  ram[14112]  = 1;
  ram[14113]  = 1;
  ram[14114]  = 1;
  ram[14115]  = 1;
  ram[14116]  = 1;
  ram[14117]  = 1;
  ram[14118]  = 1;
  ram[14119]  = 1;
  ram[14120]  = 1;
  ram[14121]  = 1;
  ram[14122]  = 1;
  ram[14123]  = 1;
  ram[14124]  = 1;
  ram[14125]  = 1;
  ram[14126]  = 1;
  ram[14127]  = 1;
  ram[14128]  = 1;
  ram[14129]  = 1;
  ram[14130]  = 1;
  ram[14131]  = 1;
  ram[14132]  = 1;
  ram[14133]  = 1;
  ram[14134]  = 1;
  ram[14135]  = 1;
  ram[14136]  = 1;
  ram[14137]  = 1;
  ram[14138]  = 1;
  ram[14139]  = 1;
  ram[14140]  = 1;
  ram[14141]  = 1;
  ram[14142]  = 1;
  ram[14143]  = 1;
  ram[14144]  = 1;
  ram[14145]  = 1;
  ram[14146]  = 1;
  ram[14147]  = 1;
  ram[14148]  = 1;
  ram[14149]  = 1;
  ram[14150]  = 1;
  ram[14151]  = 1;
  ram[14152]  = 1;
  ram[14153]  = 1;
  ram[14154]  = 1;
  ram[14155]  = 1;
  ram[14156]  = 1;
  ram[14157]  = 1;
  ram[14158]  = 1;
  ram[14159]  = 1;
  ram[14160]  = 1;
  ram[14161]  = 1;
  ram[14162]  = 1;
  ram[14163]  = 1;
  ram[14164]  = 1;
  ram[14165]  = 1;
  ram[14166]  = 1;
  ram[14167]  = 1;
  ram[14168]  = 1;
  ram[14169]  = 1;
  ram[14170]  = 1;
  ram[14171]  = 1;
  ram[14172]  = 1;
  ram[14173]  = 1;
  ram[14174]  = 1;
  ram[14175]  = 1;
  ram[14176]  = 1;
  ram[14177]  = 1;
  ram[14178]  = 1;
  ram[14179]  = 1;
  ram[14180]  = 1;
  ram[14181]  = 1;
  ram[14182]  = 1;
  ram[14183]  = 1;
  ram[14184]  = 1;
  ram[14185]  = 1;
  ram[14186]  = 1;
  ram[14187]  = 1;
  ram[14188]  = 1;
  ram[14189]  = 1;
  ram[14190]  = 1;
  ram[14191]  = 1;
  ram[14192]  = 1;
  ram[14193]  = 1;
  ram[14194]  = 1;
  ram[14195]  = 1;
  ram[14196]  = 1;
  ram[14197]  = 1;
  ram[14198]  = 1;
  ram[14199]  = 1;
  ram[14200]  = 1;
  ram[14201]  = 1;
  ram[14202]  = 1;
  ram[14203]  = 1;
  ram[14204]  = 1;
  ram[14205]  = 1;
  ram[14206]  = 1;
  ram[14207]  = 1;
  ram[14208]  = 1;
  ram[14209]  = 1;
  ram[14210]  = 1;
  ram[14211]  = 1;
  ram[14212]  = 1;
  ram[14213]  = 1;
  ram[14214]  = 1;
  ram[14215]  = 1;
  ram[14216]  = 1;
  ram[14217]  = 1;
  ram[14218]  = 1;
  ram[14219]  = 1;
  ram[14220]  = 1;
  ram[14221]  = 1;
  ram[14222]  = 1;
  ram[14223]  = 1;
  ram[14224]  = 1;
  ram[14225]  = 1;
  ram[14226]  = 1;
  ram[14227]  = 1;
  ram[14228]  = 1;
  ram[14229]  = 1;
  ram[14230]  = 1;
  ram[14231]  = 1;
  ram[14232]  = 1;
  ram[14233]  = 1;
  ram[14234]  = 1;
  ram[14235]  = 1;
  ram[14236]  = 1;
  ram[14237]  = 1;
  ram[14238]  = 1;
  ram[14239]  = 1;
  ram[14240]  = 1;
  ram[14241]  = 1;
  ram[14242]  = 1;
  ram[14243]  = 1;
  ram[14244]  = 1;
  ram[14245]  = 1;
  ram[14246]  = 1;
  ram[14247]  = 1;
  ram[14248]  = 1;
  ram[14249]  = 1;
  ram[14250]  = 1;
  ram[14251]  = 1;
  ram[14252]  = 1;
  ram[14253]  = 1;
  ram[14254]  = 1;
  ram[14255]  = 1;
  ram[14256]  = 1;
  ram[14257]  = 1;
  ram[14258]  = 1;
  ram[14259]  = 1;
  ram[14260]  = 1;
  ram[14261]  = 1;
  ram[14262]  = 1;
  ram[14263]  = 1;
  ram[14264]  = 1;
  ram[14265]  = 1;
  ram[14266]  = 1;
  ram[14267]  = 1;
  ram[14268]  = 1;
  ram[14269]  = 1;
  ram[14270]  = 1;
  ram[14271]  = 1;
  ram[14272]  = 1;
  ram[14273]  = 1;
  ram[14274]  = 1;
  ram[14275]  = 1;
  ram[14276]  = 1;
  ram[14277]  = 1;
  ram[14278]  = 1;
  ram[14279]  = 1;
  ram[14280]  = 1;
  ram[14281]  = 1;
  ram[14282]  = 1;
  ram[14283]  = 1;
  ram[14284]  = 1;
  ram[14285]  = 1;
  ram[14286]  = 1;
  ram[14287]  = 1;
  ram[14288]  = 1;
  ram[14289]  = 1;
  ram[14290]  = 1;
  ram[14291]  = 1;
  ram[14292]  = 1;
  ram[14293]  = 1;
  ram[14294]  = 1;
  ram[14295]  = 1;
  ram[14296]  = 1;
  ram[14297]  = 1;
  ram[14298]  = 1;
  ram[14299]  = 1;
  ram[14300]  = 1;
  ram[14301]  = 1;
  ram[14302]  = 1;
  ram[14303]  = 1;
  ram[14304]  = 1;
  ram[14305]  = 1;
  ram[14306]  = 1;
  ram[14307]  = 1;
  ram[14308]  = 1;
  ram[14309]  = 1;
  ram[14310]  = 1;
  ram[14311]  = 1;
  ram[14312]  = 1;
  ram[14313]  = 1;
  ram[14314]  = 1;
  ram[14315]  = 1;
  ram[14316]  = 1;
  ram[14317]  = 1;
  ram[14318]  = 1;
  ram[14319]  = 1;
  ram[14320]  = 1;
  ram[14321]  = 1;
  ram[14322]  = 1;
  ram[14323]  = 1;
  ram[14324]  = 1;
  ram[14325]  = 1;
  ram[14326]  = 1;
  ram[14327]  = 1;
  ram[14328]  = 1;
  ram[14329]  = 1;
  ram[14330]  = 1;
  ram[14331]  = 1;
  ram[14332]  = 1;
  ram[14333]  = 1;
  ram[14334]  = 1;
  ram[14335]  = 1;
  ram[14336]  = 1;
  ram[14337]  = 1;
  ram[14338]  = 1;
  ram[14339]  = 1;
  ram[14340]  = 1;
  ram[14341]  = 1;
  ram[14342]  = 1;
  ram[14343]  = 1;
  ram[14344]  = 1;
  ram[14345]  = 1;
  ram[14346]  = 1;
  ram[14347]  = 1;
  ram[14348]  = 1;
  ram[14349]  = 1;
  ram[14350]  = 1;
  ram[14351]  = 1;
  ram[14352]  = 1;
  ram[14353]  = 1;
  ram[14354]  = 1;
  ram[14355]  = 1;
  ram[14356]  = 1;
  ram[14357]  = 1;
  ram[14358]  = 1;
  ram[14359]  = 1;
  ram[14360]  = 1;
  ram[14361]  = 1;
  ram[14362]  = 1;
  ram[14363]  = 1;
  ram[14364]  = 1;
  ram[14365]  = 1;
  ram[14366]  = 1;
  ram[14367]  = 1;
  ram[14368]  = 1;
  ram[14369]  = 1;
  ram[14370]  = 1;
  ram[14371]  = 1;
  ram[14372]  = 1;
  ram[14373]  = 1;
  ram[14374]  = 1;
  ram[14375]  = 1;
  ram[14376]  = 1;
  ram[14377]  = 1;
  ram[14378]  = 1;
  ram[14379]  = 1;
  ram[14380]  = 1;
  ram[14381]  = 1;
  ram[14382]  = 1;
  ram[14383]  = 1;
  ram[14384]  = 1;
  ram[14385]  = 1;
  ram[14386]  = 1;
  ram[14387]  = 1;
  ram[14388]  = 1;
  ram[14389]  = 1;
  ram[14390]  = 1;
  ram[14391]  = 1;
  ram[14392]  = 1;
  ram[14393]  = 1;
  ram[14394]  = 1;
  ram[14395]  = 1;
  ram[14396]  = 1;
  ram[14397]  = 1;
  ram[14398]  = 1;
  ram[14399]  = 1;
  ram[14400]  = 1;
  ram[14401]  = 1;
  ram[14402]  = 1;
  ram[14403]  = 1;
  ram[14404]  = 1;
  ram[14405]  = 1;
  ram[14406]  = 1;
  ram[14407]  = 1;
  ram[14408]  = 1;
  ram[14409]  = 1;
  ram[14410]  = 1;
  ram[14411]  = 1;
  ram[14412]  = 1;
  ram[14413]  = 1;
  ram[14414]  = 1;
  ram[14415]  = 1;
  ram[14416]  = 1;
  ram[14417]  = 1;
  ram[14418]  = 1;
  ram[14419]  = 1;
  ram[14420]  = 1;
  ram[14421]  = 1;
  ram[14422]  = 1;
  ram[14423]  = 1;
  ram[14424]  = 1;
  ram[14425]  = 1;
  ram[14426]  = 1;
  ram[14427]  = 1;
  ram[14428]  = 1;
  ram[14429]  = 1;
  ram[14430]  = 1;
  ram[14431]  = 1;
  ram[14432]  = 1;
  ram[14433]  = 1;
  ram[14434]  = 1;
  ram[14435]  = 1;
  ram[14436]  = 1;
  ram[14437]  = 1;
  ram[14438]  = 1;
  ram[14439]  = 1;
  ram[14440]  = 1;
  ram[14441]  = 1;
  ram[14442]  = 1;
  ram[14443]  = 1;
  ram[14444]  = 1;
  ram[14445]  = 1;
  ram[14446]  = 1;
  ram[14447]  = 1;
  ram[14448]  = 1;
  ram[14449]  = 1;
  ram[14450]  = 1;
  ram[14451]  = 1;
  ram[14452]  = 1;
  ram[14453]  = 1;
  ram[14454]  = 1;
  ram[14455]  = 1;
  ram[14456]  = 1;
  ram[14457]  = 1;
  ram[14458]  = 1;
  ram[14459]  = 1;
  ram[14460]  = 1;
  ram[14461]  = 1;
  ram[14462]  = 1;
  ram[14463]  = 1;
  ram[14464]  = 1;
  ram[14465]  = 1;
  ram[14466]  = 1;
  ram[14467]  = 1;
  ram[14468]  = 1;
  ram[14469]  = 1;
  ram[14470]  = 1;
  ram[14471]  = 1;
  ram[14472]  = 1;
  ram[14473]  = 1;
  ram[14474]  = 1;
  ram[14475]  = 1;
  ram[14476]  = 1;
  ram[14477]  = 1;
  ram[14478]  = 1;
  ram[14479]  = 1;
  ram[14480]  = 1;
  ram[14481]  = 1;
  ram[14482]  = 1;
  ram[14483]  = 1;
  ram[14484]  = 1;
  ram[14485]  = 1;
  ram[14486]  = 1;
  ram[14487]  = 1;
  ram[14488]  = 1;
  ram[14489]  = 1;
  ram[14490]  = 1;
  ram[14491]  = 1;
  ram[14492]  = 1;
  ram[14493]  = 1;
  ram[14494]  = 1;
  ram[14495]  = 1;
  ram[14496]  = 1;
  ram[14497]  = 1;
  ram[14498]  = 1;
  ram[14499]  = 1;
  ram[14500]  = 1;
  ram[14501]  = 1;
  ram[14502]  = 1;
  ram[14503]  = 1;
  ram[14504]  = 1;
  ram[14505]  = 1;
  ram[14506]  = 1;
  ram[14507]  = 1;
  ram[14508]  = 1;
  ram[14509]  = 1;
  ram[14510]  = 1;
  ram[14511]  = 1;
  ram[14512]  = 1;
  ram[14513]  = 1;
  ram[14514]  = 1;
  ram[14515]  = 1;
  ram[14516]  = 1;
  ram[14517]  = 1;
  ram[14518]  = 1;
  ram[14519]  = 1;
  ram[14520]  = 1;
  ram[14521]  = 1;
  ram[14522]  = 1;
  ram[14523]  = 1;
  ram[14524]  = 1;
  ram[14525]  = 1;
  ram[14526]  = 1;
  ram[14527]  = 1;
  ram[14528]  = 1;
  ram[14529]  = 1;
  ram[14530]  = 1;
  ram[14531]  = 1;
  ram[14532]  = 1;
  ram[14533]  = 1;
  ram[14534]  = 1;
  ram[14535]  = 1;
  ram[14536]  = 1;
  ram[14537]  = 1;
  ram[14538]  = 1;
  ram[14539]  = 1;
  ram[14540]  = 1;
  ram[14541]  = 1;
  ram[14542]  = 1;
  ram[14543]  = 1;
  ram[14544]  = 1;
  ram[14545]  = 1;
  ram[14546]  = 1;
  ram[14547]  = 1;
  ram[14548]  = 1;
  ram[14549]  = 1;
  ram[14550]  = 1;
  ram[14551]  = 1;
  ram[14552]  = 1;
  ram[14553]  = 1;
  ram[14554]  = 1;
  ram[14555]  = 1;
  ram[14556]  = 1;
  ram[14557]  = 1;
  ram[14558]  = 1;
  ram[14559]  = 1;
  ram[14560]  = 1;
  ram[14561]  = 1;
  ram[14562]  = 1;
  ram[14563]  = 1;
  ram[14564]  = 1;
  ram[14565]  = 1;
  ram[14566]  = 1;
  ram[14567]  = 1;
  ram[14568]  = 1;
  ram[14569]  = 1;
  ram[14570]  = 1;
  ram[14571]  = 1;
  ram[14572]  = 1;
  ram[14573]  = 1;
  ram[14574]  = 1;
  ram[14575]  = 1;
  ram[14576]  = 1;
  ram[14577]  = 1;
  ram[14578]  = 1;
  ram[14579]  = 1;
  ram[14580]  = 1;
  ram[14581]  = 1;
  ram[14582]  = 1;
  ram[14583]  = 1;
  ram[14584]  = 1;
  ram[14585]  = 1;
  ram[14586]  = 1;
  ram[14587]  = 1;
  ram[14588]  = 1;
  ram[14589]  = 1;
  ram[14590]  = 1;
  ram[14591]  = 1;
  ram[14592]  = 1;
  ram[14593]  = 1;
  ram[14594]  = 1;
  ram[14595]  = 1;
  ram[14596]  = 1;
  ram[14597]  = 1;
  ram[14598]  = 1;
  ram[14599]  = 1;
  ram[14600]  = 1;
  ram[14601]  = 1;
  ram[14602]  = 1;
  ram[14603]  = 1;
  ram[14604]  = 1;
  ram[14605]  = 1;
  ram[14606]  = 1;
  ram[14607]  = 1;
  ram[14608]  = 1;
  ram[14609]  = 1;
  ram[14610]  = 1;
  ram[14611]  = 1;
  ram[14612]  = 1;
  ram[14613]  = 1;
  ram[14614]  = 1;
  ram[14615]  = 1;
  ram[14616]  = 1;
  ram[14617]  = 1;
  ram[14618]  = 1;
  ram[14619]  = 1;
  ram[14620]  = 1;
  ram[14621]  = 1;
  ram[14622]  = 1;
  ram[14623]  = 1;
  ram[14624]  = 1;
  ram[14625]  = 1;
  ram[14626]  = 1;
  ram[14627]  = 1;
  ram[14628]  = 1;
  ram[14629]  = 1;
  ram[14630]  = 1;
  ram[14631]  = 1;
  ram[14632]  = 1;
  ram[14633]  = 1;
  ram[14634]  = 1;
  ram[14635]  = 1;
  ram[14636]  = 1;
  ram[14637]  = 1;
  ram[14638]  = 1;
  ram[14639]  = 1;
  ram[14640]  = 1;
  ram[14641]  = 1;
  ram[14642]  = 1;
  ram[14643]  = 1;
  ram[14644]  = 1;
  ram[14645]  = 1;
  ram[14646]  = 1;
  ram[14647]  = 1;
  ram[14648]  = 1;
  ram[14649]  = 1;
  ram[14650]  = 1;
  ram[14651]  = 1;
  ram[14652]  = 1;
  ram[14653]  = 1;
  ram[14654]  = 1;
  ram[14655]  = 1;
  ram[14656]  = 1;
  ram[14657]  = 1;
  ram[14658]  = 1;
  ram[14659]  = 1;
  ram[14660]  = 1;
  ram[14661]  = 1;
  ram[14662]  = 1;
  ram[14663]  = 1;
  ram[14664]  = 1;
  ram[14665]  = 1;
  ram[14666]  = 1;
  ram[14667]  = 1;
  ram[14668]  = 1;
  ram[14669]  = 1;
  ram[14670]  = 1;
  ram[14671]  = 1;
  ram[14672]  = 1;
  ram[14673]  = 1;
  ram[14674]  = 1;
  ram[14675]  = 1;
  ram[14676]  = 1;
  ram[14677]  = 1;
  ram[14678]  = 1;
  ram[14679]  = 1;
  ram[14680]  = 1;
  ram[14681]  = 1;
  ram[14682]  = 1;
  ram[14683]  = 1;
  ram[14684]  = 1;
  ram[14685]  = 1;
  ram[14686]  = 1;
  ram[14687]  = 1;
  ram[14688]  = 1;
  ram[14689]  = 1;
  ram[14690]  = 1;
  ram[14691]  = 1;
  ram[14692]  = 1;
  ram[14693]  = 1;
  ram[14694]  = 1;
  ram[14695]  = 1;
  ram[14696]  = 1;
  ram[14697]  = 1;
  ram[14698]  = 1;
  ram[14699]  = 1;
  ram[14700]  = 1;
  ram[14701]  = 1;
  ram[14702]  = 1;
  ram[14703]  = 1;
  ram[14704]  = 1;
  ram[14705]  = 1;
  ram[14706]  = 1;
  ram[14707]  = 1;
  ram[14708]  = 1;
  ram[14709]  = 1;
  ram[14710]  = 1;
  ram[14711]  = 1;
  ram[14712]  = 1;
  ram[14713]  = 1;
  ram[14714]  = 1;
  ram[14715]  = 1;
  ram[14716]  = 1;
  ram[14717]  = 1;
  ram[14718]  = 1;
  ram[14719]  = 1;
  ram[14720]  = 1;
  ram[14721]  = 1;
  ram[14722]  = 1;
  ram[14723]  = 1;
  ram[14724]  = 1;
  ram[14725]  = 1;
  ram[14726]  = 1;
  ram[14727]  = 1;
  ram[14728]  = 1;
  ram[14729]  = 1;
  ram[14730]  = 1;
  ram[14731]  = 1;
  ram[14732]  = 1;
  ram[14733]  = 1;
  ram[14734]  = 1;
  ram[14735]  = 1;
  ram[14736]  = 1;
  ram[14737]  = 1;
  ram[14738]  = 1;
  ram[14739]  = 1;
  ram[14740]  = 1;
  ram[14741]  = 1;
  ram[14742]  = 1;
  ram[14743]  = 1;
  ram[14744]  = 1;
  ram[14745]  = 1;
  ram[14746]  = 1;
  ram[14747]  = 1;
  ram[14748]  = 1;
  ram[14749]  = 1;
  ram[14750]  = 1;
  ram[14751]  = 1;
  ram[14752]  = 1;
  ram[14753]  = 1;
  ram[14754]  = 1;
  ram[14755]  = 1;
  ram[14756]  = 1;
  ram[14757]  = 1;
  ram[14758]  = 1;
  ram[14759]  = 1;
  ram[14760]  = 1;
  ram[14761]  = 1;
  ram[14762]  = 1;
  ram[14763]  = 1;
  ram[14764]  = 1;
  ram[14765]  = 1;
  ram[14766]  = 1;
  ram[14767]  = 1;
  ram[14768]  = 1;
  ram[14769]  = 1;
  ram[14770]  = 1;
  ram[14771]  = 1;
  ram[14772]  = 1;
  ram[14773]  = 1;
  ram[14774]  = 1;
  ram[14775]  = 1;
  ram[14776]  = 1;
  ram[14777]  = 1;
  ram[14778]  = 1;
  ram[14779]  = 1;
  ram[14780]  = 1;
  ram[14781]  = 1;
  ram[14782]  = 1;
  ram[14783]  = 1;
  ram[14784]  = 1;
  ram[14785]  = 1;
  ram[14786]  = 1;
  ram[14787]  = 1;
  ram[14788]  = 1;
  ram[14789]  = 1;
  ram[14790]  = 1;
  ram[14791]  = 1;
  ram[14792]  = 1;
  ram[14793]  = 1;
  ram[14794]  = 1;
  ram[14795]  = 1;
  ram[14796]  = 1;
  ram[14797]  = 1;
  ram[14798]  = 1;
  ram[14799]  = 1;
  ram[14800]  = 1;
  ram[14801]  = 1;
  ram[14802]  = 1;
  ram[14803]  = 1;
  ram[14804]  = 1;
  ram[14805]  = 1;
  ram[14806]  = 1;
  ram[14807]  = 1;
  ram[14808]  = 1;
  ram[14809]  = 1;
  ram[14810]  = 1;
  ram[14811]  = 1;
  ram[14812]  = 1;
  ram[14813]  = 1;
  ram[14814]  = 1;
  ram[14815]  = 1;
  ram[14816]  = 1;
  ram[14817]  = 1;
  ram[14818]  = 1;
  ram[14819]  = 1;
  ram[14820]  = 1;
  ram[14821]  = 1;
  ram[14822]  = 1;
  ram[14823]  = 1;
  ram[14824]  = 1;
  ram[14825]  = 1;
  ram[14826]  = 1;
  ram[14827]  = 1;
  ram[14828]  = 1;
  ram[14829]  = 1;
  ram[14830]  = 1;
  ram[14831]  = 1;
  ram[14832]  = 1;
  ram[14833]  = 1;
  ram[14834]  = 1;
  ram[14835]  = 1;
  ram[14836]  = 1;
  ram[14837]  = 1;
  ram[14838]  = 1;
  ram[14839]  = 1;
  ram[14840]  = 1;
  ram[14841]  = 1;
  ram[14842]  = 1;
  ram[14843]  = 1;
  ram[14844]  = 1;
  ram[14845]  = 1;
  ram[14846]  = 1;
  ram[14847]  = 1;
  ram[14848]  = 1;
  ram[14849]  = 1;
  ram[14850]  = 1;
  ram[14851]  = 1;
  ram[14852]  = 1;
  ram[14853]  = 1;
  ram[14854]  = 1;
  ram[14855]  = 1;
  ram[14856]  = 1;
  ram[14857]  = 1;
  ram[14858]  = 1;
  ram[14859]  = 1;
  ram[14860]  = 1;
  ram[14861]  = 1;
  ram[14862]  = 1;
  ram[14863]  = 1;
  ram[14864]  = 1;
  ram[14865]  = 1;
  ram[14866]  = 1;
  ram[14867]  = 1;
  ram[14868]  = 1;
  ram[14869]  = 1;
  ram[14870]  = 1;
  ram[14871]  = 1;
  ram[14872]  = 1;
  ram[14873]  = 1;
  ram[14874]  = 1;
  ram[14875]  = 1;
  ram[14876]  = 1;
  ram[14877]  = 1;
  ram[14878]  = 1;
  ram[14879]  = 1;
  ram[14880]  = 1;
  ram[14881]  = 1;
  ram[14882]  = 1;
  ram[14883]  = 1;
  ram[14884]  = 1;
  ram[14885]  = 1;
  ram[14886]  = 1;
  ram[14887]  = 1;
  ram[14888]  = 1;
  ram[14889]  = 1;
  ram[14890]  = 1;
  ram[14891]  = 1;
  ram[14892]  = 1;
  ram[14893]  = 1;
  ram[14894]  = 1;
  ram[14895]  = 1;
  ram[14896]  = 1;
  ram[14897]  = 1;
  ram[14898]  = 1;
  ram[14899]  = 1;
  ram[14900]  = 1;
  ram[14901]  = 1;
  ram[14902]  = 1;
  ram[14903]  = 1;
  ram[14904]  = 1;
  ram[14905]  = 1;
  ram[14906]  = 1;
  ram[14907]  = 1;
  ram[14908]  = 1;
  ram[14909]  = 1;
  ram[14910]  = 1;
  ram[14911]  = 1;
  ram[14912]  = 1;
  ram[14913]  = 1;
  ram[14914]  = 1;
  ram[14915]  = 1;
  ram[14916]  = 1;
  ram[14917]  = 1;
  ram[14918]  = 1;
  ram[14919]  = 1;
  ram[14920]  = 1;
  ram[14921]  = 1;
  ram[14922]  = 1;
  ram[14923]  = 1;
  ram[14924]  = 1;
  ram[14925]  = 1;
  ram[14926]  = 1;
  ram[14927]  = 1;
  ram[14928]  = 1;
  ram[14929]  = 1;
  ram[14930]  = 1;
  ram[14931]  = 1;
  ram[14932]  = 1;
  ram[14933]  = 1;
  ram[14934]  = 1;
  ram[14935]  = 1;
  ram[14936]  = 1;
  ram[14937]  = 1;
  ram[14938]  = 1;
  ram[14939]  = 1;
  ram[14940]  = 1;
  ram[14941]  = 1;
  ram[14942]  = 1;
  ram[14943]  = 1;
  ram[14944]  = 1;
  ram[14945]  = 1;
  ram[14946]  = 1;
  ram[14947]  = 1;
  ram[14948]  = 1;
  ram[14949]  = 1;
  ram[14950]  = 1;
  ram[14951]  = 1;
  ram[14952]  = 1;
  ram[14953]  = 1;
  ram[14954]  = 1;
  ram[14955]  = 1;
  ram[14956]  = 1;
  ram[14957]  = 1;
  ram[14958]  = 1;
  ram[14959]  = 1;
  ram[14960]  = 1;
  ram[14961]  = 1;
  ram[14962]  = 1;
  ram[14963]  = 1;
  ram[14964]  = 1;
  ram[14965]  = 1;
  ram[14966]  = 1;
  ram[14967]  = 1;
  ram[14968]  = 1;
  ram[14969]  = 1;
  ram[14970]  = 1;
  ram[14971]  = 1;
  ram[14972]  = 1;
  ram[14973]  = 1;
  ram[14974]  = 1;
  ram[14975]  = 1;
  ram[14976]  = 1;
  ram[14977]  = 1;
  ram[14978]  = 1;
  ram[14979]  = 1;
  ram[14980]  = 1;
  ram[14981]  = 1;
  ram[14982]  = 1;
  ram[14983]  = 1;
  ram[14984]  = 1;
  ram[14985]  = 1;
  ram[14986]  = 1;
  ram[14987]  = 1;
  ram[14988]  = 1;
  ram[14989]  = 1;
  ram[14990]  = 1;
  ram[14991]  = 1;
  ram[14992]  = 1;
  ram[14993]  = 1;
  ram[14994]  = 1;
  ram[14995]  = 1;
  ram[14996]  = 1;
  ram[14997]  = 1;
  ram[14998]  = 1;
  ram[14999]  = 1;
  ram[15000]  = 1;
  ram[15001]  = 1;
  ram[15002]  = 1;
  ram[15003]  = 1;
  ram[15004]  = 1;
  ram[15005]  = 1;
  ram[15006]  = 1;
  ram[15007]  = 1;
  ram[15008]  = 1;
  ram[15009]  = 1;
  ram[15010]  = 1;
  ram[15011]  = 1;
  ram[15012]  = 1;
  ram[15013]  = 1;
  ram[15014]  = 1;
  ram[15015]  = 1;
  ram[15016]  = 1;
  ram[15017]  = 1;
  ram[15018]  = 1;
  ram[15019]  = 1;
  ram[15020]  = 1;
  ram[15021]  = 1;
  ram[15022]  = 1;
  ram[15023]  = 1;
  ram[15024]  = 1;
  ram[15025]  = 1;
  ram[15026]  = 1;
  ram[15027]  = 1;
  ram[15028]  = 1;
  ram[15029]  = 1;
  ram[15030]  = 1;
  ram[15031]  = 1;
  ram[15032]  = 1;
  ram[15033]  = 1;
  ram[15034]  = 1;
  ram[15035]  = 1;
  ram[15036]  = 1;
  ram[15037]  = 1;
  ram[15038]  = 1;
  ram[15039]  = 1;
  ram[15040]  = 1;
  ram[15041]  = 1;
  ram[15042]  = 1;
  ram[15043]  = 1;
  ram[15044]  = 1;
  ram[15045]  = 1;
  ram[15046]  = 1;
  ram[15047]  = 1;
  ram[15048]  = 1;
  ram[15049]  = 1;
  ram[15050]  = 1;
  ram[15051]  = 1;
  ram[15052]  = 1;
  ram[15053]  = 1;
  ram[15054]  = 1;
  ram[15055]  = 1;
  ram[15056]  = 1;
  ram[15057]  = 1;
  ram[15058]  = 1;
  ram[15059]  = 1;
  ram[15060]  = 1;
  ram[15061]  = 1;
  ram[15062]  = 1;
  ram[15063]  = 1;
  ram[15064]  = 1;
  ram[15065]  = 1;
  ram[15066]  = 1;
  ram[15067]  = 1;
  ram[15068]  = 1;
  ram[15069]  = 1;
  ram[15070]  = 1;
  ram[15071]  = 1;
  ram[15072]  = 1;
  ram[15073]  = 1;
  ram[15074]  = 1;
  ram[15075]  = 1;
  ram[15076]  = 1;
  ram[15077]  = 1;
  ram[15078]  = 1;
  ram[15079]  = 1;
  ram[15080]  = 1;
  ram[15081]  = 1;
  ram[15082]  = 1;
  ram[15083]  = 1;
  ram[15084]  = 1;
  ram[15085]  = 1;
  ram[15086]  = 1;
  ram[15087]  = 1;
  ram[15088]  = 1;
  ram[15089]  = 1;
  ram[15090]  = 1;
  ram[15091]  = 1;
  ram[15092]  = 1;
  ram[15093]  = 1;
  ram[15094]  = 1;
  ram[15095]  = 1;
  ram[15096]  = 1;
  ram[15097]  = 1;
  ram[15098]  = 1;
  ram[15099]  = 1;
  ram[15100]  = 1;
  ram[15101]  = 1;
  ram[15102]  = 1;
  ram[15103]  = 1;
  ram[15104]  = 1;
  ram[15105]  = 1;
  ram[15106]  = 1;
  ram[15107]  = 1;
  ram[15108]  = 1;
  ram[15109]  = 1;
  ram[15110]  = 1;
  ram[15111]  = 1;
  ram[15112]  = 1;
  ram[15113]  = 1;
  ram[15114]  = 1;
  ram[15115]  = 1;
  ram[15116]  = 1;
  ram[15117]  = 1;
  ram[15118]  = 1;
  ram[15119]  = 1;
  ram[15120]  = 1;
  ram[15121]  = 1;
  ram[15122]  = 1;
  ram[15123]  = 1;
  ram[15124]  = 1;
  ram[15125]  = 1;
  ram[15126]  = 1;
  ram[15127]  = 1;
  ram[15128]  = 1;
  ram[15129]  = 1;
  ram[15130]  = 1;
  ram[15131]  = 1;
  ram[15132]  = 1;
  ram[15133]  = 1;
  ram[15134]  = 1;
  ram[15135]  = 1;
  ram[15136]  = 1;
  ram[15137]  = 1;
  ram[15138]  = 1;
  ram[15139]  = 1;
  ram[15140]  = 1;
  ram[15141]  = 1;
  ram[15142]  = 1;
  ram[15143]  = 1;
  ram[15144]  = 1;
  ram[15145]  = 1;
  ram[15146]  = 1;
  ram[15147]  = 1;
  ram[15148]  = 1;
  ram[15149]  = 1;
  ram[15150]  = 1;
  ram[15151]  = 1;
  ram[15152]  = 1;
  ram[15153]  = 1;
  ram[15154]  = 1;
  ram[15155]  = 1;
  ram[15156]  = 1;
  ram[15157]  = 1;
  ram[15158]  = 1;
  ram[15159]  = 1;
  ram[15160]  = 1;
  ram[15161]  = 1;
  ram[15162]  = 1;
  ram[15163]  = 1;
  ram[15164]  = 1;
  ram[15165]  = 1;
  ram[15166]  = 1;
  ram[15167]  = 1;
  ram[15168]  = 1;
  ram[15169]  = 1;
  ram[15170]  = 1;
  ram[15171]  = 1;
  ram[15172]  = 1;
  ram[15173]  = 1;
  ram[15174]  = 1;
  ram[15175]  = 1;
  ram[15176]  = 1;
  ram[15177]  = 1;
  ram[15178]  = 1;
  ram[15179]  = 1;
  ram[15180]  = 1;
  ram[15181]  = 1;
  ram[15182]  = 1;
  ram[15183]  = 1;
  ram[15184]  = 1;
  ram[15185]  = 1;
  ram[15186]  = 1;
  ram[15187]  = 1;
  ram[15188]  = 1;
  ram[15189]  = 1;
  ram[15190]  = 1;
  ram[15191]  = 1;
  ram[15192]  = 1;
  ram[15193]  = 1;
  ram[15194]  = 1;
  ram[15195]  = 1;
  ram[15196]  = 1;
  ram[15197]  = 1;
  ram[15198]  = 1;
  ram[15199]  = 1;
  ram[15200]  = 1;
  ram[15201]  = 1;
  ram[15202]  = 1;
  ram[15203]  = 1;
  ram[15204]  = 1;
  ram[15205]  = 1;
  ram[15206]  = 1;
  ram[15207]  = 1;
  ram[15208]  = 1;
  ram[15209]  = 1;
  ram[15210]  = 1;
  ram[15211]  = 1;
  ram[15212]  = 1;
  ram[15213]  = 1;
  ram[15214]  = 1;
  ram[15215]  = 1;
  ram[15216]  = 1;
  ram[15217]  = 1;
  ram[15218]  = 1;
  ram[15219]  = 1;
  ram[15220]  = 1;
  ram[15221]  = 1;
  ram[15222]  = 1;
  ram[15223]  = 1;
  ram[15224]  = 1;
  ram[15225]  = 1;
  ram[15226]  = 1;
  ram[15227]  = 1;
  ram[15228]  = 1;
  ram[15229]  = 1;
  ram[15230]  = 1;
  ram[15231]  = 1;
  ram[15232]  = 1;
  ram[15233]  = 1;
  ram[15234]  = 1;
  ram[15235]  = 1;
  ram[15236]  = 1;
  ram[15237]  = 1;
  ram[15238]  = 1;
  ram[15239]  = 1;
  ram[15240]  = 1;
  ram[15241]  = 1;
  ram[15242]  = 1;
  ram[15243]  = 1;
  ram[15244]  = 1;
  ram[15245]  = 1;
  ram[15246]  = 1;
  ram[15247]  = 1;
  ram[15248]  = 1;
  ram[15249]  = 1;
  ram[15250]  = 1;
  ram[15251]  = 1;
  ram[15252]  = 1;
  ram[15253]  = 1;
  ram[15254]  = 1;
  ram[15255]  = 1;
  ram[15256]  = 1;
  ram[15257]  = 1;
  ram[15258]  = 1;
  ram[15259]  = 1;
  ram[15260]  = 1;
  ram[15261]  = 1;
  ram[15262]  = 1;
  ram[15263]  = 1;
  ram[15264]  = 1;
  ram[15265]  = 1;
  ram[15266]  = 1;
  ram[15267]  = 1;
  ram[15268]  = 1;
  ram[15269]  = 1;
  ram[15270]  = 1;
  ram[15271]  = 1;
  ram[15272]  = 1;
  ram[15273]  = 1;
  ram[15274]  = 1;
  ram[15275]  = 1;
  ram[15276]  = 1;
  ram[15277]  = 1;
  ram[15278]  = 1;
  ram[15279]  = 1;
  ram[15280]  = 1;
  ram[15281]  = 1;
  ram[15282]  = 1;
  ram[15283]  = 1;
  ram[15284]  = 1;
  ram[15285]  = 1;
  ram[15286]  = 1;
  ram[15287]  = 1;
  ram[15288]  = 1;
  ram[15289]  = 1;
  ram[15290]  = 1;
  ram[15291]  = 1;
  ram[15292]  = 1;
  ram[15293]  = 1;
  ram[15294]  = 1;
  ram[15295]  = 1;
  ram[15296]  = 1;
  ram[15297]  = 1;
  ram[15298]  = 1;
  ram[15299]  = 1;
  ram[15300]  = 1;
  ram[15301]  = 1;
  ram[15302]  = 1;
  ram[15303]  = 1;
  ram[15304]  = 1;
  ram[15305]  = 1;
  ram[15306]  = 1;
  ram[15307]  = 1;
  ram[15308]  = 1;
  ram[15309]  = 1;
  ram[15310]  = 1;
  ram[15311]  = 1;
  ram[15312]  = 1;
  ram[15313]  = 1;
  ram[15314]  = 1;
  ram[15315]  = 1;
  ram[15316]  = 1;
  ram[15317]  = 1;
  ram[15318]  = 1;
  ram[15319]  = 1;
  ram[15320]  = 1;
  ram[15321]  = 1;
  ram[15322]  = 1;
  ram[15323]  = 1;
  ram[15324]  = 1;
  ram[15325]  = 1;
  ram[15326]  = 1;
  ram[15327]  = 1;
  ram[15328]  = 1;
  ram[15329]  = 1;
  ram[15330]  = 1;
  ram[15331]  = 1;
  ram[15332]  = 1;
  ram[15333]  = 1;
  ram[15334]  = 1;
  ram[15335]  = 1;
  ram[15336]  = 1;
  ram[15337]  = 1;
  ram[15338]  = 1;
  ram[15339]  = 1;
  ram[15340]  = 1;
  ram[15341]  = 1;
  ram[15342]  = 1;
  ram[15343]  = 1;
  ram[15344]  = 1;
  ram[15345]  = 1;
  ram[15346]  = 1;
  ram[15347]  = 1;
  ram[15348]  = 1;
  ram[15349]  = 1;
  ram[15350]  = 1;
  ram[15351]  = 1;
  ram[15352]  = 1;
  ram[15353]  = 1;
  ram[15354]  = 1;
  ram[15355]  = 1;
  ram[15356]  = 1;
  ram[15357]  = 1;
  ram[15358]  = 1;
  ram[15359]  = 1;
  ram[15360]  = 1;
  ram[15361]  = 1;
  ram[15362]  = 1;
  ram[15363]  = 1;
  ram[15364]  = 1;
  ram[15365]  = 1;
  ram[15366]  = 1;
  ram[15367]  = 1;
  ram[15368]  = 1;
  ram[15369]  = 1;
  ram[15370]  = 1;
  ram[15371]  = 1;
  ram[15372]  = 1;
  ram[15373]  = 1;
  ram[15374]  = 1;
  ram[15375]  = 1;
  ram[15376]  = 1;
  ram[15377]  = 1;
  ram[15378]  = 1;
  ram[15379]  = 1;
  ram[15380]  = 1;
  ram[15381]  = 1;
  ram[15382]  = 1;
  ram[15383]  = 1;
  ram[15384]  = 1;
  ram[15385]  = 1;
  ram[15386]  = 1;
  ram[15387]  = 1;
  ram[15388]  = 1;
  ram[15389]  = 1;
  ram[15390]  = 1;
  ram[15391]  = 1;
  ram[15392]  = 1;
  ram[15393]  = 1;
  ram[15394]  = 1;
  ram[15395]  = 1;
  ram[15396]  = 1;
  ram[15397]  = 1;
  ram[15398]  = 1;
  ram[15399]  = 1;
  ram[15400]  = 1;
  ram[15401]  = 1;
  ram[15402]  = 1;
  ram[15403]  = 1;
  ram[15404]  = 1;
  ram[15405]  = 1;
  ram[15406]  = 1;
  ram[15407]  = 1;
  ram[15408]  = 1;
  ram[15409]  = 1;
  ram[15410]  = 1;
  ram[15411]  = 1;
  ram[15412]  = 1;
  ram[15413]  = 1;
  ram[15414]  = 1;
  ram[15415]  = 1;
  ram[15416]  = 1;
  ram[15417]  = 1;
  ram[15418]  = 1;
  ram[15419]  = 1;
  ram[15420]  = 1;
  ram[15421]  = 1;
  ram[15422]  = 1;
  ram[15423]  = 1;
  ram[15424]  = 1;
  ram[15425]  = 1;
  ram[15426]  = 1;
  ram[15427]  = 1;
  ram[15428]  = 1;
  ram[15429]  = 1;
  ram[15430]  = 1;
  ram[15431]  = 1;
  ram[15432]  = 1;
  ram[15433]  = 1;
  ram[15434]  = 1;
  ram[15435]  = 1;
  ram[15436]  = 1;
  ram[15437]  = 1;
  ram[15438]  = 1;
  ram[15439]  = 1;
  ram[15440]  = 1;
  ram[15441]  = 1;
  ram[15442]  = 1;
  ram[15443]  = 1;
  ram[15444]  = 1;
  ram[15445]  = 1;
  ram[15446]  = 1;
  ram[15447]  = 1;
  ram[15448]  = 1;
  ram[15449]  = 1;
  ram[15450]  = 1;
  ram[15451]  = 1;
  ram[15452]  = 1;
  ram[15453]  = 1;
  ram[15454]  = 1;
  ram[15455]  = 1;
  ram[15456]  = 1;
  ram[15457]  = 1;
  ram[15458]  = 1;
  ram[15459]  = 1;
  ram[15460]  = 1;
  ram[15461]  = 1;
  ram[15462]  = 1;
  ram[15463]  = 1;
  ram[15464]  = 1;
  ram[15465]  = 1;
  ram[15466]  = 1;
  ram[15467]  = 1;
  ram[15468]  = 1;
  ram[15469]  = 1;
  ram[15470]  = 1;
  ram[15471]  = 1;
  ram[15472]  = 1;
  ram[15473]  = 1;
  ram[15474]  = 1;
  ram[15475]  = 1;
  ram[15476]  = 1;
  ram[15477]  = 1;
  ram[15478]  = 1;
  ram[15479]  = 1;
  ram[15480]  = 1;
  ram[15481]  = 1;
  ram[15482]  = 1;
  ram[15483]  = 1;
  ram[15484]  = 1;
  ram[15485]  = 1;
  ram[15486]  = 1;
  ram[15487]  = 1;
  ram[15488]  = 1;
  ram[15489]  = 1;
  ram[15490]  = 1;
  ram[15491]  = 1;
  ram[15492]  = 1;
  ram[15493]  = 1;
  ram[15494]  = 1;
  ram[15495]  = 1;
  ram[15496]  = 1;
  ram[15497]  = 1;
  ram[15498]  = 1;
  ram[15499]  = 1;
  ram[15500]  = 1;
  ram[15501]  = 1;
  ram[15502]  = 1;
  ram[15503]  = 1;
  ram[15504]  = 1;
  ram[15505]  = 1;
  ram[15506]  = 1;
  ram[15507]  = 1;
  ram[15508]  = 1;
  ram[15509]  = 1;
  ram[15510]  = 1;
  ram[15511]  = 1;
  ram[15512]  = 1;
  ram[15513]  = 1;
  ram[15514]  = 1;
  ram[15515]  = 1;
  ram[15516]  = 1;
  ram[15517]  = 1;
  ram[15518]  = 1;
  ram[15519]  = 1;
  ram[15520]  = 1;
  ram[15521]  = 1;
  ram[15522]  = 1;
  ram[15523]  = 1;
  ram[15524]  = 1;
  ram[15525]  = 1;
  ram[15526]  = 1;
  ram[15527]  = 1;
  ram[15528]  = 1;
  ram[15529]  = 1;
  ram[15530]  = 1;
  ram[15531]  = 1;
  ram[15532]  = 1;
  ram[15533]  = 1;
  ram[15534]  = 1;
  ram[15535]  = 1;
  ram[15536]  = 1;
  ram[15537]  = 1;
  ram[15538]  = 1;
  ram[15539]  = 1;
  ram[15540]  = 1;
  ram[15541]  = 1;
  ram[15542]  = 1;
  ram[15543]  = 1;
  ram[15544]  = 1;
  ram[15545]  = 1;
  ram[15546]  = 1;
  ram[15547]  = 1;
  ram[15548]  = 1;
  ram[15549]  = 1;
  ram[15550]  = 1;
  ram[15551]  = 1;
  ram[15552]  = 1;
  ram[15553]  = 1;
  ram[15554]  = 1;
  ram[15555]  = 1;
  ram[15556]  = 1;
  ram[15557]  = 1;
  ram[15558]  = 1;
  ram[15559]  = 1;
  ram[15560]  = 1;
  ram[15561]  = 1;
  ram[15562]  = 1;
  ram[15563]  = 1;
  ram[15564]  = 1;
  ram[15565]  = 1;
  ram[15566]  = 1;
  ram[15567]  = 1;
  ram[15568]  = 1;
  ram[15569]  = 1;
  ram[15570]  = 1;
  ram[15571]  = 1;
  ram[15572]  = 1;
  ram[15573]  = 1;
  ram[15574]  = 1;
  ram[15575]  = 1;
  ram[15576]  = 1;
  ram[15577]  = 1;
  ram[15578]  = 1;
  ram[15579]  = 1;
  ram[15580]  = 1;
  ram[15581]  = 1;
  ram[15582]  = 1;
  ram[15583]  = 1;
  ram[15584]  = 1;
  ram[15585]  = 1;
  ram[15586]  = 1;
  ram[15587]  = 1;
  ram[15588]  = 1;
  ram[15589]  = 1;
  ram[15590]  = 1;
  ram[15591]  = 1;
  ram[15592]  = 1;
  ram[15593]  = 1;
  ram[15594]  = 1;
  ram[15595]  = 1;
  ram[15596]  = 1;
  ram[15597]  = 1;
  ram[15598]  = 1;
  ram[15599]  = 1;
  ram[15600]  = 1;
  ram[15601]  = 1;
  ram[15602]  = 1;
  ram[15603]  = 1;
  ram[15604]  = 1;
  ram[15605]  = 1;
  ram[15606]  = 1;
  ram[15607]  = 1;
  ram[15608]  = 1;
  ram[15609]  = 1;
  ram[15610]  = 1;
  ram[15611]  = 1;
  ram[15612]  = 1;
  ram[15613]  = 1;
  ram[15614]  = 1;
  ram[15615]  = 1;
  ram[15616]  = 1;
  ram[15617]  = 1;
  ram[15618]  = 1;
  ram[15619]  = 1;
  ram[15620]  = 1;
  ram[15621]  = 1;
  ram[15622]  = 1;
  ram[15623]  = 1;
  ram[15624]  = 1;
  ram[15625]  = 1;
  ram[15626]  = 1;
  ram[15627]  = 1;
  ram[15628]  = 1;
  ram[15629]  = 1;
  ram[15630]  = 1;
  ram[15631]  = 1;
  ram[15632]  = 1;
  ram[15633]  = 1;
  ram[15634]  = 1;
  ram[15635]  = 1;
  ram[15636]  = 1;
  ram[15637]  = 1;
  ram[15638]  = 1;
  ram[15639]  = 1;
  ram[15640]  = 1;
  ram[15641]  = 1;
  ram[15642]  = 1;
  ram[15643]  = 1;
  ram[15644]  = 1;
  ram[15645]  = 1;
  ram[15646]  = 1;
  ram[15647]  = 1;
  ram[15648]  = 1;
  ram[15649]  = 1;
  ram[15650]  = 1;
  ram[15651]  = 1;
  ram[15652]  = 1;
  ram[15653]  = 1;
  ram[15654]  = 1;
  ram[15655]  = 1;
  ram[15656]  = 1;
  ram[15657]  = 1;
  ram[15658]  = 1;
  ram[15659]  = 1;
  ram[15660]  = 1;
  ram[15661]  = 1;
  ram[15662]  = 1;
  ram[15663]  = 1;
  ram[15664]  = 1;
  ram[15665]  = 1;
  ram[15666]  = 1;
  ram[15667]  = 1;
  ram[15668]  = 1;
  ram[15669]  = 1;
  ram[15670]  = 1;
  ram[15671]  = 1;
  ram[15672]  = 1;
  ram[15673]  = 1;
  ram[15674]  = 1;
  ram[15675]  = 1;
  ram[15676]  = 1;
  ram[15677]  = 1;
  ram[15678]  = 1;
  ram[15679]  = 1;
  ram[15680]  = 1;
  ram[15681]  = 1;
  ram[15682]  = 1;
  ram[15683]  = 1;
  ram[15684]  = 1;
  ram[15685]  = 1;
  ram[15686]  = 1;
  ram[15687]  = 1;
  ram[15688]  = 1;
  ram[15689]  = 1;
  ram[15690]  = 1;
  ram[15691]  = 1;
  ram[15692]  = 1;
  ram[15693]  = 1;
  ram[15694]  = 1;
  ram[15695]  = 1;
  ram[15696]  = 1;
  ram[15697]  = 1;
  ram[15698]  = 1;
  ram[15699]  = 1;
  ram[15700]  = 1;
  ram[15701]  = 1;
  ram[15702]  = 1;
  ram[15703]  = 1;
  ram[15704]  = 1;
  ram[15705]  = 1;
  ram[15706]  = 1;
  ram[15707]  = 1;
  ram[15708]  = 1;
  ram[15709]  = 1;
  ram[15710]  = 1;
  ram[15711]  = 1;
  ram[15712]  = 1;
  ram[15713]  = 1;
  ram[15714]  = 1;
  ram[15715]  = 1;
  ram[15716]  = 1;
  ram[15717]  = 1;
  ram[15718]  = 1;
  ram[15719]  = 1;
  ram[15720]  = 1;
  ram[15721]  = 1;
  ram[15722]  = 1;
  ram[15723]  = 1;
  ram[15724]  = 1;
  ram[15725]  = 1;
  ram[15726]  = 1;
  ram[15727]  = 1;
  ram[15728]  = 1;
  ram[15729]  = 1;
  ram[15730]  = 1;
  ram[15731]  = 1;
  ram[15732]  = 1;
  ram[15733]  = 1;
  ram[15734]  = 1;
  ram[15735]  = 1;
  ram[15736]  = 1;
  ram[15737]  = 1;
  ram[15738]  = 1;
  ram[15739]  = 1;
  ram[15740]  = 1;
  ram[15741]  = 1;
  ram[15742]  = 1;
  ram[15743]  = 1;
  ram[15744]  = 1;
  ram[15745]  = 1;
  ram[15746]  = 1;
  ram[15747]  = 1;
  ram[15748]  = 1;
  ram[15749]  = 1;
  ram[15750]  = 1;
  ram[15751]  = 1;
  ram[15752]  = 1;
  ram[15753]  = 1;
  ram[15754]  = 1;
  ram[15755]  = 1;
  ram[15756]  = 1;
  ram[15757]  = 1;
  ram[15758]  = 1;
  ram[15759]  = 1;
  ram[15760]  = 1;
  ram[15761]  = 1;
  ram[15762]  = 1;
  ram[15763]  = 1;
  ram[15764]  = 1;
  ram[15765]  = 1;
  ram[15766]  = 1;
  ram[15767]  = 1;
  ram[15768]  = 1;
  ram[15769]  = 1;
  ram[15770]  = 1;
  ram[15771]  = 1;
  ram[15772]  = 1;
  ram[15773]  = 1;
  ram[15774]  = 1;
  ram[15775]  = 1;
  ram[15776]  = 1;
  ram[15777]  = 1;
  ram[15778]  = 1;
  ram[15779]  = 1;
  ram[15780]  = 1;
  ram[15781]  = 1;
  ram[15782]  = 1;
  ram[15783]  = 1;
  ram[15784]  = 1;
  ram[15785]  = 1;
  ram[15786]  = 1;
  ram[15787]  = 1;
  ram[15788]  = 1;
  ram[15789]  = 1;
  ram[15790]  = 1;
  ram[15791]  = 1;
  ram[15792]  = 1;
  ram[15793]  = 1;
  ram[15794]  = 1;
  ram[15795]  = 1;
  ram[15796]  = 1;
  ram[15797]  = 1;
  ram[15798]  = 1;
  ram[15799]  = 1;
  ram[15800]  = 1;
  ram[15801]  = 1;
  ram[15802]  = 1;
  ram[15803]  = 1;
  ram[15804]  = 1;
  ram[15805]  = 1;
  ram[15806]  = 1;
  ram[15807]  = 1;
  ram[15808]  = 1;
  ram[15809]  = 1;
  ram[15810]  = 1;
  ram[15811]  = 1;
  ram[15812]  = 1;
  ram[15813]  = 1;
  ram[15814]  = 1;
  ram[15815]  = 1;
  ram[15816]  = 1;
  ram[15817]  = 1;
  ram[15818]  = 1;
  ram[15819]  = 1;
  ram[15820]  = 1;
  ram[15821]  = 1;
  ram[15822]  = 1;
  ram[15823]  = 1;
  ram[15824]  = 1;
  ram[15825]  = 1;
  ram[15826]  = 1;
  ram[15827]  = 1;
  ram[15828]  = 1;
  ram[15829]  = 1;
  ram[15830]  = 1;
  ram[15831]  = 1;
  ram[15832]  = 1;
  ram[15833]  = 1;
  ram[15834]  = 1;
  ram[15835]  = 1;
  ram[15836]  = 1;
  ram[15837]  = 1;
  ram[15838]  = 1;
  ram[15839]  = 1;
  ram[15840]  = 1;
  ram[15841]  = 1;
  ram[15842]  = 1;
  ram[15843]  = 1;
  ram[15844]  = 1;
  ram[15845]  = 1;
  ram[15846]  = 1;
  ram[15847]  = 1;
  ram[15848]  = 1;
  ram[15849]  = 1;
  ram[15850]  = 1;
  ram[15851]  = 1;
  ram[15852]  = 1;
  ram[15853]  = 1;
  ram[15854]  = 1;
  ram[15855]  = 1;
  ram[15856]  = 1;
  ram[15857]  = 1;
  ram[15858]  = 1;
  ram[15859]  = 1;
  ram[15860]  = 1;
  ram[15861]  = 1;
  ram[15862]  = 1;
  ram[15863]  = 1;
  ram[15864]  = 1;
  ram[15865]  = 1;
  ram[15866]  = 1;
  ram[15867]  = 1;
  ram[15868]  = 1;
  ram[15869]  = 1;
  ram[15870]  = 1;
  ram[15871]  = 1;
  ram[15872]  = 1;
  ram[15873]  = 1;
  ram[15874]  = 1;
  ram[15875]  = 1;
  ram[15876]  = 1;
  ram[15877]  = 1;
  ram[15878]  = 1;
  ram[15879]  = 1;
  ram[15880]  = 1;
  ram[15881]  = 1;
  ram[15882]  = 1;
  ram[15883]  = 1;
  ram[15884]  = 1;
  ram[15885]  = 1;
  ram[15886]  = 1;
  ram[15887]  = 1;
  ram[15888]  = 1;
  ram[15889]  = 1;
  ram[15890]  = 1;
  ram[15891]  = 1;
  ram[15892]  = 1;
  ram[15893]  = 1;
  ram[15894]  = 1;
  ram[15895]  = 1;
  ram[15896]  = 1;
  ram[15897]  = 1;
  ram[15898]  = 1;
  ram[15899]  = 1;
  ram[15900]  = 1;
  ram[15901]  = 1;
  ram[15902]  = 1;
  ram[15903]  = 1;
  ram[15904]  = 1;
  ram[15905]  = 1;
  ram[15906]  = 1;
  ram[15907]  = 1;
  ram[15908]  = 1;
  ram[15909]  = 1;
  ram[15910]  = 1;
  ram[15911]  = 1;
  ram[15912]  = 1;
  ram[15913]  = 1;
  ram[15914]  = 1;
  ram[15915]  = 1;
  ram[15916]  = 1;
  ram[15917]  = 1;
  ram[15918]  = 1;
  ram[15919]  = 1;
  ram[15920]  = 1;
  ram[15921]  = 1;
  ram[15922]  = 1;
  ram[15923]  = 1;
  ram[15924]  = 1;
  ram[15925]  = 1;
  ram[15926]  = 1;
  ram[15927]  = 1;
  ram[15928]  = 1;
  ram[15929]  = 1;
  ram[15930]  = 1;
  ram[15931]  = 1;
  ram[15932]  = 1;
  ram[15933]  = 1;
  ram[15934]  = 1;
  ram[15935]  = 1;
  ram[15936]  = 1;
  ram[15937]  = 1;
  ram[15938]  = 1;
  ram[15939]  = 1;
  ram[15940]  = 1;
  ram[15941]  = 1;
  ram[15942]  = 1;
  ram[15943]  = 1;
  ram[15944]  = 1;
  ram[15945]  = 1;
  ram[15946]  = 1;
  ram[15947]  = 1;
  ram[15948]  = 1;
  ram[15949]  = 1;
  ram[15950]  = 1;
  ram[15951]  = 1;
  ram[15952]  = 1;
  ram[15953]  = 1;
  ram[15954]  = 1;
  ram[15955]  = 1;
  ram[15956]  = 1;
  ram[15957]  = 1;
  ram[15958]  = 1;
  ram[15959]  = 1;
  ram[15960]  = 1;
  ram[15961]  = 1;
  ram[15962]  = 1;
  ram[15963]  = 1;
  ram[15964]  = 1;
  ram[15965]  = 1;
  ram[15966]  = 1;
  ram[15967]  = 1;
  ram[15968]  = 1;
  ram[15969]  = 1;
  ram[15970]  = 1;
  ram[15971]  = 1;
  ram[15972]  = 1;
  ram[15973]  = 1;
  ram[15974]  = 1;
  ram[15975]  = 1;
  ram[15976]  = 1;
  ram[15977]  = 1;
  ram[15978]  = 1;
  ram[15979]  = 1;
  ram[15980]  = 1;
  ram[15981]  = 1;
  ram[15982]  = 1;
  ram[15983]  = 1;
  ram[15984]  = 1;
  ram[15985]  = 1;
  ram[15986]  = 1;
  ram[15987]  = 1;
  ram[15988]  = 1;
  ram[15989]  = 1;
  ram[15990]  = 1;
  ram[15991]  = 1;
  ram[15992]  = 1;
  ram[15993]  = 1;
  ram[15994]  = 1;
  ram[15995]  = 1;
  ram[15996]  = 1;
  ram[15997]  = 1;
  ram[15998]  = 1;
  ram[15999]  = 1;
  ram[16000]  = 1;
  ram[16001]  = 1;
  ram[16002]  = 1;
  ram[16003]  = 1;
  ram[16004]  = 1;
  ram[16005]  = 1;
  ram[16006]  = 1;
  ram[16007]  = 1;
  ram[16008]  = 1;
  ram[16009]  = 1;
  ram[16010]  = 1;
  ram[16011]  = 1;
  ram[16012]  = 1;
  ram[16013]  = 1;
  ram[16014]  = 1;
  ram[16015]  = 1;
  ram[16016]  = 1;
  ram[16017]  = 1;
  ram[16018]  = 1;
  ram[16019]  = 1;
  ram[16020]  = 1;
  ram[16021]  = 1;
  ram[16022]  = 1;
  ram[16023]  = 1;
  ram[16024]  = 1;
  ram[16025]  = 1;
  ram[16026]  = 1;
  ram[16027]  = 1;
  ram[16028]  = 1;
  ram[16029]  = 1;
  ram[16030]  = 1;
  ram[16031]  = 1;
  ram[16032]  = 1;
  ram[16033]  = 1;
  ram[16034]  = 1;
  ram[16035]  = 1;
  ram[16036]  = 1;
  ram[16037]  = 1;
  ram[16038]  = 1;
  ram[16039]  = 1;
  ram[16040]  = 1;
  ram[16041]  = 1;
  ram[16042]  = 1;
  ram[16043]  = 1;
  ram[16044]  = 1;
  ram[16045]  = 1;
  ram[16046]  = 1;
  ram[16047]  = 1;
  ram[16048]  = 1;
  ram[16049]  = 1;
  ram[16050]  = 1;
  ram[16051]  = 1;
  ram[16052]  = 1;
  ram[16053]  = 1;
  ram[16054]  = 1;
  ram[16055]  = 1;
  ram[16056]  = 1;
  ram[16057]  = 1;
  ram[16058]  = 1;
  ram[16059]  = 1;
  ram[16060]  = 1;
  ram[16061]  = 1;
  ram[16062]  = 1;
  ram[16063]  = 1;
  ram[16064]  = 1;
  ram[16065]  = 1;
  ram[16066]  = 1;
  ram[16067]  = 1;
  ram[16068]  = 1;
  ram[16069]  = 1;
  ram[16070]  = 1;
  ram[16071]  = 1;
  ram[16072]  = 1;
  ram[16073]  = 1;
  ram[16074]  = 1;
  ram[16075]  = 1;
  ram[16076]  = 1;
  ram[16077]  = 1;
  ram[16078]  = 1;
  ram[16079]  = 1;
  ram[16080]  = 1;
  ram[16081]  = 1;
  ram[16082]  = 1;
  ram[16083]  = 1;
  ram[16084]  = 1;
  ram[16085]  = 1;
  ram[16086]  = 1;
  ram[16087]  = 1;
  ram[16088]  = 1;
  ram[16089]  = 1;
  ram[16090]  = 1;
  ram[16091]  = 1;
  ram[16092]  = 1;
  ram[16093]  = 1;
  ram[16094]  = 1;
  ram[16095]  = 1;
  ram[16096]  = 1;
  ram[16097]  = 1;
  ram[16098]  = 1;
  ram[16099]  = 1;
  ram[16100]  = 1;
  ram[16101]  = 1;
  ram[16102]  = 1;
  ram[16103]  = 1;
  ram[16104]  = 1;
  ram[16105]  = 1;
  ram[16106]  = 1;
  ram[16107]  = 1;
  ram[16108]  = 1;
  ram[16109]  = 1;
  ram[16110]  = 1;
  ram[16111]  = 1;
  ram[16112]  = 1;
  ram[16113]  = 1;
  ram[16114]  = 1;
  ram[16115]  = 1;
  ram[16116]  = 1;
  ram[16117]  = 1;
  ram[16118]  = 1;
  ram[16119]  = 1;
  ram[16120]  = 1;
  ram[16121]  = 1;
  ram[16122]  = 1;
  ram[16123]  = 1;
  ram[16124]  = 1;
  ram[16125]  = 1;
  ram[16126]  = 1;
  ram[16127]  = 1;
  ram[16128]  = 1;
  ram[16129]  = 1;
  ram[16130]  = 1;
  ram[16131]  = 1;
  ram[16132]  = 1;
  ram[16133]  = 1;
  ram[16134]  = 1;
  ram[16135]  = 1;
  ram[16136]  = 1;
  ram[16137]  = 1;
  ram[16138]  = 1;
  ram[16139]  = 1;
  ram[16140]  = 1;
  ram[16141]  = 1;
  ram[16142]  = 1;
  ram[16143]  = 1;
  ram[16144]  = 1;
  ram[16145]  = 1;
  ram[16146]  = 1;
  ram[16147]  = 1;
  ram[16148]  = 1;
  ram[16149]  = 1;
  ram[16150]  = 1;
  ram[16151]  = 1;
  ram[16152]  = 1;
  ram[16153]  = 1;
  ram[16154]  = 1;
  ram[16155]  = 1;
  ram[16156]  = 1;
  ram[16157]  = 1;
  ram[16158]  = 1;
  ram[16159]  = 1;
  ram[16160]  = 1;
  ram[16161]  = 1;
  ram[16162]  = 1;
  ram[16163]  = 1;
  ram[16164]  = 1;
  ram[16165]  = 1;
  ram[16166]  = 1;
  ram[16167]  = 1;
  ram[16168]  = 1;
  ram[16169]  = 1;
  ram[16170]  = 1;
  ram[16171]  = 1;
  ram[16172]  = 1;
  ram[16173]  = 1;
  ram[16174]  = 1;
  ram[16175]  = 1;
  ram[16176]  = 1;
  ram[16177]  = 1;
  ram[16178]  = 1;
  ram[16179]  = 1;
  ram[16180]  = 1;
  ram[16181]  = 1;
  ram[16182]  = 1;
  ram[16183]  = 1;
  ram[16184]  = 1;
  ram[16185]  = 1;
  ram[16186]  = 1;
  ram[16187]  = 1;
  ram[16188]  = 1;
  ram[16189]  = 1;
  ram[16190]  = 1;
  ram[16191]  = 1;
  ram[16192]  = 1;
  ram[16193]  = 1;
  ram[16194]  = 1;
  ram[16195]  = 1;
  ram[16196]  = 1;
  ram[16197]  = 1;
  ram[16198]  = 1;
  ram[16199]  = 1;
  ram[16200]  = 1;
  ram[16201]  = 1;
  ram[16202]  = 1;
  ram[16203]  = 1;
  ram[16204]  = 1;
  ram[16205]  = 1;
  ram[16206]  = 1;
  ram[16207]  = 1;
  ram[16208]  = 1;
  ram[16209]  = 1;
  ram[16210]  = 1;
  ram[16211]  = 1;
  ram[16212]  = 1;
  ram[16213]  = 1;
  ram[16214]  = 1;
  ram[16215]  = 1;
  ram[16216]  = 1;
  ram[16217]  = 1;
  ram[16218]  = 1;
  ram[16219]  = 1;
  ram[16220]  = 1;
  ram[16221]  = 1;
  ram[16222]  = 1;
  ram[16223]  = 1;
  ram[16224]  = 1;
  ram[16225]  = 1;
  ram[16226]  = 1;
  ram[16227]  = 1;
  ram[16228]  = 1;
  ram[16229]  = 1;
  ram[16230]  = 1;
  ram[16231]  = 1;
  ram[16232]  = 1;
  ram[16233]  = 1;
  ram[16234]  = 1;
  ram[16235]  = 1;
  ram[16236]  = 1;
  ram[16237]  = 1;
  ram[16238]  = 1;
  ram[16239]  = 1;
  ram[16240]  = 1;
  ram[16241]  = 1;
  ram[16242]  = 1;
  ram[16243]  = 1;
  ram[16244]  = 1;
  ram[16245]  = 1;
  ram[16246]  = 1;
  ram[16247]  = 1;
  ram[16248]  = 1;
  ram[16249]  = 1;
  ram[16250]  = 1;
  ram[16251]  = 1;
  ram[16252]  = 1;
  ram[16253]  = 1;
  ram[16254]  = 1;
  ram[16255]  = 1;
  ram[16256]  = 1;
  ram[16257]  = 1;
  ram[16258]  = 1;
  ram[16259]  = 1;
  ram[16260]  = 1;
  ram[16261]  = 1;
  ram[16262]  = 1;
  ram[16263]  = 1;
  ram[16264]  = 1;
  ram[16265]  = 1;
  ram[16266]  = 1;
  ram[16267]  = 1;
  ram[16268]  = 1;
  ram[16269]  = 1;
  ram[16270]  = 1;
  ram[16271]  = 1;
  ram[16272]  = 1;
  ram[16273]  = 1;
  ram[16274]  = 1;
  ram[16275]  = 1;
  ram[16276]  = 1;
  ram[16277]  = 1;
  ram[16278]  = 1;
  ram[16279]  = 1;
  ram[16280]  = 1;
  ram[16281]  = 1;
  ram[16282]  = 1;
  ram[16283]  = 1;
  ram[16284]  = 1;
  ram[16285]  = 1;
  ram[16286]  = 1;
  ram[16287]  = 1;
  ram[16288]  = 1;
  ram[16289]  = 1;
  ram[16290]  = 1;
  ram[16291]  = 1;
  ram[16292]  = 1;
  ram[16293]  = 1;
  ram[16294]  = 1;
  ram[16295]  = 1;
  ram[16296]  = 1;
  ram[16297]  = 1;
  ram[16298]  = 1;
  ram[16299]  = 1;
  ram[16300]  = 1;
  ram[16301]  = 1;
  ram[16302]  = 1;
  ram[16303]  = 1;
  ram[16304]  = 1;
  ram[16305]  = 1;
  ram[16306]  = 1;
  ram[16307]  = 1;
  ram[16308]  = 1;
  ram[16309]  = 1;
  ram[16310]  = 1;
  ram[16311]  = 1;
  ram[16312]  = 1;
  ram[16313]  = 1;
  ram[16314]  = 1;
  ram[16315]  = 1;
  ram[16316]  = 1;
  ram[16317]  = 1;
  ram[16318]  = 1;
  ram[16319]  = 1;
  ram[16320]  = 1;
  ram[16321]  = 1;
  ram[16322]  = 1;
  ram[16323]  = 1;
  ram[16324]  = 1;
  ram[16325]  = 1;
  ram[16326]  = 1;
  ram[16327]  = 1;
  ram[16328]  = 1;
  ram[16329]  = 1;
  ram[16330]  = 1;
  ram[16331]  = 1;
  ram[16332]  = 1;
  ram[16333]  = 1;
  ram[16334]  = 1;
  ram[16335]  = 1;
  ram[16336]  = 1;
  ram[16337]  = 1;
  ram[16338]  = 1;
  ram[16339]  = 1;
  ram[16340]  = 1;
  ram[16341]  = 1;
  ram[16342]  = 1;
  ram[16343]  = 1;
  ram[16344]  = 1;
  ram[16345]  = 1;
  ram[16346]  = 1;
  ram[16347]  = 1;
  ram[16348]  = 1;
  ram[16349]  = 1;
  ram[16350]  = 1;
  ram[16351]  = 1;
  ram[16352]  = 1;
  ram[16353]  = 1;
  ram[16354]  = 1;
  ram[16355]  = 1;
  ram[16356]  = 1;
  ram[16357]  = 1;
  ram[16358]  = 1;
  ram[16359]  = 1;
  ram[16360]  = 1;
  ram[16361]  = 1;
  ram[16362]  = 1;
  ram[16363]  = 1;
  ram[16364]  = 1;
  ram[16365]  = 1;
  ram[16366]  = 1;
  ram[16367]  = 1;
  ram[16368]  = 1;
  ram[16369]  = 1;
  ram[16370]  = 1;
  ram[16371]  = 1;
  ram[16372]  = 1;
  ram[16373]  = 1;
  ram[16374]  = 1;
  ram[16375]  = 1;
  ram[16376]  = 1;
  ram[16377]  = 1;
  ram[16378]  = 1;
  ram[16379]  = 1;
  ram[16380]  = 1;
  ram[16381]  = 1;
  ram[16382]  = 1;
  ram[16383]  = 1;
  ram[16384]  = 1;
  ram[16385]  = 1;
  ram[16386]  = 1;
  ram[16387]  = 1;
  ram[16388]  = 1;
  ram[16389]  = 1;
  ram[16390]  = 1;
  ram[16391]  = 1;
  ram[16392]  = 1;
  ram[16393]  = 1;
  ram[16394]  = 1;
  ram[16395]  = 1;
  ram[16396]  = 1;
  ram[16397]  = 1;
  ram[16398]  = 1;
  ram[16399]  = 1;
  ram[16400]  = 1;
  ram[16401]  = 1;
  ram[16402]  = 1;
  ram[16403]  = 1;
  ram[16404]  = 1;
  ram[16405]  = 1;
  ram[16406]  = 1;
  ram[16407]  = 1;
  ram[16408]  = 1;
  ram[16409]  = 1;
  ram[16410]  = 1;
  ram[16411]  = 1;
  ram[16412]  = 1;
  ram[16413]  = 1;
  ram[16414]  = 1;
  ram[16415]  = 1;
  ram[16416]  = 1;
  ram[16417]  = 1;
  ram[16418]  = 1;
  ram[16419]  = 1;
  ram[16420]  = 1;
  ram[16421]  = 1;
  ram[16422]  = 1;
  ram[16423]  = 1;
  ram[16424]  = 1;
  ram[16425]  = 1;
  ram[16426]  = 1;
  ram[16427]  = 1;
  ram[16428]  = 1;
  ram[16429]  = 1;
  ram[16430]  = 1;
  ram[16431]  = 1;
  ram[16432]  = 1;
  ram[16433]  = 1;
  ram[16434]  = 1;
  ram[16435]  = 1;
  ram[16436]  = 1;
  ram[16437]  = 1;
  ram[16438]  = 1;
  ram[16439]  = 1;
  ram[16440]  = 1;
  ram[16441]  = 1;
  ram[16442]  = 1;
  ram[16443]  = 1;
  ram[16444]  = 1;
  ram[16445]  = 1;
  ram[16446]  = 1;
  ram[16447]  = 1;
  ram[16448]  = 1;
  ram[16449]  = 1;
  ram[16450]  = 1;
  ram[16451]  = 1;
  ram[16452]  = 1;
  ram[16453]  = 1;
  ram[16454]  = 1;
  ram[16455]  = 1;
  ram[16456]  = 1;
  ram[16457]  = 1;
  ram[16458]  = 1;
  ram[16459]  = 1;
  ram[16460]  = 1;
  ram[16461]  = 1;
  ram[16462]  = 1;
  ram[16463]  = 1;
  ram[16464]  = 1;
  ram[16465]  = 1;
  ram[16466]  = 1;
  ram[16467]  = 1;
  ram[16468]  = 1;
  ram[16469]  = 1;
  ram[16470]  = 1;
  ram[16471]  = 1;
  ram[16472]  = 1;
  ram[16473]  = 1;
  ram[16474]  = 1;
  ram[16475]  = 1;
  ram[16476]  = 1;
  ram[16477]  = 1;
  ram[16478]  = 1;
  ram[16479]  = 1;
  ram[16480]  = 1;
  ram[16481]  = 1;
  ram[16482]  = 1;
  ram[16483]  = 1;
  ram[16484]  = 1;
  ram[16485]  = 1;
  ram[16486]  = 1;
  ram[16487]  = 1;
  ram[16488]  = 1;
  ram[16489]  = 1;
  ram[16490]  = 1;
  ram[16491]  = 1;
  ram[16492]  = 1;
  ram[16493]  = 1;
  ram[16494]  = 1;
  ram[16495]  = 1;
  ram[16496]  = 1;
  ram[16497]  = 1;
  ram[16498]  = 1;
  ram[16499]  = 1;
  ram[16500]  = 1;
  ram[16501]  = 1;
  ram[16502]  = 1;
  ram[16503]  = 1;
  ram[16504]  = 1;
  ram[16505]  = 1;
  ram[16506]  = 1;
  ram[16507]  = 1;
  ram[16508]  = 1;
  ram[16509]  = 1;
  ram[16510]  = 1;
  ram[16511]  = 1;
  ram[16512]  = 1;
  ram[16513]  = 1;
  ram[16514]  = 1;
  ram[16515]  = 1;
  ram[16516]  = 1;
  ram[16517]  = 1;
  ram[16518]  = 1;
  ram[16519]  = 1;
  ram[16520]  = 1;
  ram[16521]  = 1;
  ram[16522]  = 1;
  ram[16523]  = 1;
  ram[16524]  = 1;
  ram[16525]  = 1;
  ram[16526]  = 1;
  ram[16527]  = 1;
  ram[16528]  = 1;
  ram[16529]  = 1;
  ram[16530]  = 1;
  ram[16531]  = 1;
  ram[16532]  = 1;
  ram[16533]  = 1;
  ram[16534]  = 1;
  ram[16535]  = 1;
  ram[16536]  = 1;
  ram[16537]  = 1;
  ram[16538]  = 1;
  ram[16539]  = 1;
  ram[16540]  = 1;
  ram[16541]  = 1;
  ram[16542]  = 1;
  ram[16543]  = 1;
  ram[16544]  = 1;
  ram[16545]  = 1;
  ram[16546]  = 1;
  ram[16547]  = 1;
  ram[16548]  = 1;
  ram[16549]  = 1;
  ram[16550]  = 1;
  ram[16551]  = 1;
  ram[16552]  = 1;
  ram[16553]  = 1;
  ram[16554]  = 1;
  ram[16555]  = 1;
  ram[16556]  = 1;
  ram[16557]  = 1;
  ram[16558]  = 1;
  ram[16559]  = 1;
  ram[16560]  = 1;
  ram[16561]  = 1;
  ram[16562]  = 1;
  ram[16563]  = 1;
  ram[16564]  = 1;
  ram[16565]  = 1;
  ram[16566]  = 1;
  ram[16567]  = 1;
  ram[16568]  = 1;
  ram[16569]  = 1;
  ram[16570]  = 1;
  ram[16571]  = 1;
  ram[16572]  = 1;
  ram[16573]  = 1;
  ram[16574]  = 1;
  ram[16575]  = 1;
  ram[16576]  = 1;
  ram[16577]  = 1;
  ram[16578]  = 1;
  ram[16579]  = 1;
  ram[16580]  = 1;
  ram[16581]  = 1;
  ram[16582]  = 1;
  ram[16583]  = 1;
  ram[16584]  = 1;
  ram[16585]  = 1;
  ram[16586]  = 1;
  ram[16587]  = 1;
  ram[16588]  = 1;
  ram[16589]  = 1;
  ram[16590]  = 1;
  ram[16591]  = 1;
  ram[16592]  = 1;
  ram[16593]  = 1;
  ram[16594]  = 1;
  ram[16595]  = 1;
  ram[16596]  = 1;
  ram[16597]  = 1;
  ram[16598]  = 1;
  ram[16599]  = 1;
  ram[16600]  = 1;
  ram[16601]  = 1;
  ram[16602]  = 1;
  ram[16603]  = 1;
  ram[16604]  = 1;
  ram[16605]  = 1;
  ram[16606]  = 1;
  ram[16607]  = 1;
  ram[16608]  = 1;
  ram[16609]  = 1;
  ram[16610]  = 1;
  ram[16611]  = 1;
  ram[16612]  = 1;
  ram[16613]  = 1;
  ram[16614]  = 1;
  ram[16615]  = 1;
  ram[16616]  = 1;
  ram[16617]  = 1;
  ram[16618]  = 1;
  ram[16619]  = 1;
  ram[16620]  = 1;
  ram[16621]  = 1;
  ram[16622]  = 1;
  ram[16623]  = 1;
  ram[16624]  = 1;
  ram[16625]  = 1;
  ram[16626]  = 1;
  ram[16627]  = 1;
  ram[16628]  = 1;
  ram[16629]  = 1;
  ram[16630]  = 1;
  ram[16631]  = 1;
  ram[16632]  = 1;
  ram[16633]  = 1;
  ram[16634]  = 1;
  ram[16635]  = 1;
  ram[16636]  = 1;
  ram[16637]  = 1;
  ram[16638]  = 1;
  ram[16639]  = 1;
  ram[16640]  = 1;
  ram[16641]  = 1;
  ram[16642]  = 1;
  ram[16643]  = 1;
  ram[16644]  = 1;
  ram[16645]  = 1;
  ram[16646]  = 1;
  ram[16647]  = 1;
  ram[16648]  = 1;
  ram[16649]  = 1;
  ram[16650]  = 1;
  ram[16651]  = 1;
  ram[16652]  = 1;
  ram[16653]  = 1;
  ram[16654]  = 1;
  ram[16655]  = 1;
  ram[16656]  = 1;
  ram[16657]  = 1;
  ram[16658]  = 1;
  ram[16659]  = 1;
  ram[16660]  = 1;
  ram[16661]  = 1;
  ram[16662]  = 1;
  ram[16663]  = 1;
  ram[16664]  = 1;
  ram[16665]  = 1;
  ram[16666]  = 1;
  ram[16667]  = 1;
  ram[16668]  = 1;
  ram[16669]  = 1;
  ram[16670]  = 1;
  ram[16671]  = 1;
  ram[16672]  = 1;
  ram[16673]  = 1;
  ram[16674]  = 1;
  ram[16675]  = 1;
  ram[16676]  = 1;
  ram[16677]  = 1;
  ram[16678]  = 1;
  ram[16679]  = 1;
  ram[16680]  = 1;
  ram[16681]  = 1;
  ram[16682]  = 1;
  ram[16683]  = 1;
  ram[16684]  = 1;
  ram[16685]  = 1;
  ram[16686]  = 1;
  ram[16687]  = 1;
  ram[16688]  = 1;
  ram[16689]  = 1;
  ram[16690]  = 1;
  ram[16691]  = 1;
  ram[16692]  = 1;
  ram[16693]  = 1;
  ram[16694]  = 1;
  ram[16695]  = 1;
  ram[16696]  = 1;
  ram[16697]  = 1;
  ram[16698]  = 1;
  ram[16699]  = 1;
  ram[16700]  = 1;
  ram[16701]  = 1;
  ram[16702]  = 1;
  ram[16703]  = 1;
  ram[16704]  = 1;
  ram[16705]  = 1;
  ram[16706]  = 1;
  ram[16707]  = 1;
  ram[16708]  = 1;
  ram[16709]  = 1;
  ram[16710]  = 1;
  ram[16711]  = 1;
  ram[16712]  = 1;
  ram[16713]  = 1;
  ram[16714]  = 1;
  ram[16715]  = 1;
  ram[16716]  = 1;
  ram[16717]  = 1;
  ram[16718]  = 1;
  ram[16719]  = 1;
  ram[16720]  = 1;
  ram[16721]  = 1;
  ram[16722]  = 1;
  ram[16723]  = 1;
  ram[16724]  = 1;
  ram[16725]  = 1;
  ram[16726]  = 1;
  ram[16727]  = 1;
  ram[16728]  = 1;
  ram[16729]  = 1;
  ram[16730]  = 1;
  ram[16731]  = 1;
  ram[16732]  = 1;
  ram[16733]  = 1;
  ram[16734]  = 1;
  ram[16735]  = 1;
  ram[16736]  = 1;
  ram[16737]  = 1;
  ram[16738]  = 1;
  ram[16739]  = 1;
  ram[16740]  = 1;
  ram[16741]  = 1;
  ram[16742]  = 1;
  ram[16743]  = 1;
  ram[16744]  = 1;
  ram[16745]  = 1;
  ram[16746]  = 1;
  ram[16747]  = 1;
  ram[16748]  = 1;
  ram[16749]  = 1;
  ram[16750]  = 1;
  ram[16751]  = 1;
  ram[16752]  = 1;
  ram[16753]  = 1;
  ram[16754]  = 1;
  ram[16755]  = 1;
  ram[16756]  = 1;
  ram[16757]  = 1;
  ram[16758]  = 1;
  ram[16759]  = 1;
  ram[16760]  = 1;
  ram[16761]  = 1;
  ram[16762]  = 1;
  ram[16763]  = 1;
  ram[16764]  = 1;
  ram[16765]  = 1;
  ram[16766]  = 1;
  ram[16767]  = 1;
  ram[16768]  = 1;
  ram[16769]  = 1;
  ram[16770]  = 1;
  ram[16771]  = 1;
  ram[16772]  = 1;
  ram[16773]  = 1;
  ram[16774]  = 1;
  ram[16775]  = 1;
  ram[16776]  = 1;
  ram[16777]  = 1;
  ram[16778]  = 1;
  ram[16779]  = 1;
  ram[16780]  = 1;
  ram[16781]  = 1;
  ram[16782]  = 1;
  ram[16783]  = 1;
  ram[16784]  = 1;
  ram[16785]  = 1;
  ram[16786]  = 1;
  ram[16787]  = 1;
  ram[16788]  = 1;
  ram[16789]  = 1;
  ram[16790]  = 1;
  ram[16791]  = 1;
  ram[16792]  = 1;
  ram[16793]  = 1;
  ram[16794]  = 1;
  ram[16795]  = 1;
  ram[16796]  = 1;
  ram[16797]  = 1;
  ram[16798]  = 1;
  ram[16799]  = 1;
  ram[16800]  = 1;
  ram[16801]  = 1;
  ram[16802]  = 1;
  ram[16803]  = 1;
  ram[16804]  = 1;
  ram[16805]  = 1;
  ram[16806]  = 1;
  ram[16807]  = 1;
  ram[16808]  = 1;
  ram[16809]  = 1;
  ram[16810]  = 1;
  ram[16811]  = 1;
  ram[16812]  = 1;
  ram[16813]  = 1;
  ram[16814]  = 1;
  ram[16815]  = 1;
  ram[16816]  = 1;
  ram[16817]  = 1;
  ram[16818]  = 1;
  ram[16819]  = 1;
  ram[16820]  = 1;
  ram[16821]  = 1;
  ram[16822]  = 1;
  ram[16823]  = 1;
  ram[16824]  = 1;
  ram[16825]  = 1;
  ram[16826]  = 1;
  ram[16827]  = 1;
  ram[16828]  = 1;
  ram[16829]  = 1;
  ram[16830]  = 1;
  ram[16831]  = 1;
  ram[16832]  = 1;
  ram[16833]  = 1;
  ram[16834]  = 1;
  ram[16835]  = 1;
  ram[16836]  = 1;
  ram[16837]  = 1;
  ram[16838]  = 1;
  ram[16839]  = 1;
  ram[16840]  = 1;
  ram[16841]  = 1;
  ram[16842]  = 1;
  ram[16843]  = 1;
  ram[16844]  = 1;
  ram[16845]  = 1;
  ram[16846]  = 1;
  ram[16847]  = 1;
  ram[16848]  = 1;
  ram[16849]  = 1;
  ram[16850]  = 1;
  ram[16851]  = 1;
  ram[16852]  = 1;
  ram[16853]  = 1;
  ram[16854]  = 1;
  ram[16855]  = 1;
  ram[16856]  = 1;
  ram[16857]  = 1;
  ram[16858]  = 1;
  ram[16859]  = 1;
  ram[16860]  = 1;
  ram[16861]  = 1;
  ram[16862]  = 1;
  ram[16863]  = 1;
  ram[16864]  = 1;
  ram[16865]  = 1;
  ram[16866]  = 1;
  ram[16867]  = 1;
  ram[16868]  = 1;
  ram[16869]  = 1;
  ram[16870]  = 1;
  ram[16871]  = 1;
  ram[16872]  = 1;
  ram[16873]  = 1;
  ram[16874]  = 1;
  ram[16875]  = 1;
  ram[16876]  = 1;
  ram[16877]  = 1;
  ram[16878]  = 1;
  ram[16879]  = 1;
  ram[16880]  = 1;
  ram[16881]  = 1;
  ram[16882]  = 1;
  ram[16883]  = 1;
  ram[16884]  = 1;
  ram[16885]  = 1;
  ram[16886]  = 1;
  ram[16887]  = 1;
  ram[16888]  = 1;
  ram[16889]  = 1;
  ram[16890]  = 1;
  ram[16891]  = 1;
  ram[16892]  = 1;
  ram[16893]  = 1;
  ram[16894]  = 1;
  ram[16895]  = 1;
  ram[16896]  = 1;
  ram[16897]  = 1;
  ram[16898]  = 1;
  ram[16899]  = 1;
  ram[16900]  = 1;
  ram[16901]  = 1;
  ram[16902]  = 1;
  ram[16903]  = 1;
  ram[16904]  = 1;
  ram[16905]  = 1;
  ram[16906]  = 1;
  ram[16907]  = 1;
  ram[16908]  = 1;
  ram[16909]  = 1;
  ram[16910]  = 1;
  ram[16911]  = 1;
  ram[16912]  = 1;
  ram[16913]  = 1;
  ram[16914]  = 1;
  ram[16915]  = 1;
  ram[16916]  = 1;
  ram[16917]  = 1;
  ram[16918]  = 1;
  ram[16919]  = 1;
  ram[16920]  = 1;
  ram[16921]  = 1;
  ram[16922]  = 1;
  ram[16923]  = 1;
  ram[16924]  = 1;
  ram[16925]  = 1;
  ram[16926]  = 1;
  ram[16927]  = 1;
  ram[16928]  = 1;
  ram[16929]  = 1;
  ram[16930]  = 1;
  ram[16931]  = 1;
  ram[16932]  = 1;
  ram[16933]  = 1;
  ram[16934]  = 1;
  ram[16935]  = 1;
  ram[16936]  = 1;
  ram[16937]  = 1;
  ram[16938]  = 1;
  ram[16939]  = 1;
  ram[16940]  = 1;
  ram[16941]  = 1;
  ram[16942]  = 1;
  ram[16943]  = 1;
  ram[16944]  = 1;
  ram[16945]  = 1;
  ram[16946]  = 1;
  ram[16947]  = 1;
  ram[16948]  = 1;
  ram[16949]  = 1;
  ram[16950]  = 1;
  ram[16951]  = 1;
  ram[16952]  = 1;
  ram[16953]  = 1;
  ram[16954]  = 1;
  ram[16955]  = 1;
  ram[16956]  = 1;
  ram[16957]  = 1;
  ram[16958]  = 1;
  ram[16959]  = 1;
  ram[16960]  = 1;
  ram[16961]  = 1;
  ram[16962]  = 1;
  ram[16963]  = 1;
  ram[16964]  = 1;
  ram[16965]  = 1;
  ram[16966]  = 1;
  ram[16967]  = 1;
  ram[16968]  = 1;
  ram[16969]  = 1;
  ram[16970]  = 1;
  ram[16971]  = 1;
  ram[16972]  = 1;
  ram[16973]  = 1;
  ram[16974]  = 1;
  ram[16975]  = 1;
  ram[16976]  = 1;
  ram[16977]  = 1;
  ram[16978]  = 1;
  ram[16979]  = 1;
  ram[16980]  = 1;
  ram[16981]  = 1;
  ram[16982]  = 1;
  ram[16983]  = 1;
  ram[16984]  = 1;
  ram[16985]  = 1;
  ram[16986]  = 1;
  ram[16987]  = 1;
  ram[16988]  = 1;
  ram[16989]  = 1;
  ram[16990]  = 1;
  ram[16991]  = 1;
  ram[16992]  = 1;
  ram[16993]  = 1;
  ram[16994]  = 1;
  ram[16995]  = 1;
  ram[16996]  = 1;
  ram[16997]  = 1;
  ram[16998]  = 1;
  ram[16999]  = 1;
  ram[17000]  = 1;
  ram[17001]  = 1;
  ram[17002]  = 1;
  ram[17003]  = 1;
  ram[17004]  = 1;
  ram[17005]  = 1;
  ram[17006]  = 1;
  ram[17007]  = 1;
  ram[17008]  = 1;
  ram[17009]  = 1;
  ram[17010]  = 1;
  ram[17011]  = 1;
  ram[17012]  = 1;
  ram[17013]  = 1;
  ram[17014]  = 1;
  ram[17015]  = 1;
  ram[17016]  = 1;
  ram[17017]  = 1;
  ram[17018]  = 1;
  ram[17019]  = 1;
  ram[17020]  = 1;
  ram[17021]  = 1;
  ram[17022]  = 1;
  ram[17023]  = 1;
  ram[17024]  = 1;
  ram[17025]  = 1;
  ram[17026]  = 1;
  ram[17027]  = 1;
  ram[17028]  = 1;
  ram[17029]  = 1;
  ram[17030]  = 1;
  ram[17031]  = 1;
  ram[17032]  = 1;
  ram[17033]  = 1;
  ram[17034]  = 1;
  ram[17035]  = 1;
  ram[17036]  = 1;
  ram[17037]  = 1;
  ram[17038]  = 1;
  ram[17039]  = 1;
  ram[17040]  = 1;
  ram[17041]  = 1;
  ram[17042]  = 1;
  ram[17043]  = 1;
  ram[17044]  = 1;
  ram[17045]  = 1;
  ram[17046]  = 1;
  ram[17047]  = 1;
  ram[17048]  = 1;
  ram[17049]  = 1;
  ram[17050]  = 1;
  ram[17051]  = 1;
  ram[17052]  = 1;
  ram[17053]  = 1;
  ram[17054]  = 1;
  ram[17055]  = 1;
  ram[17056]  = 1;
  ram[17057]  = 1;
  ram[17058]  = 1;
  ram[17059]  = 1;
  ram[17060]  = 1;
  ram[17061]  = 1;
  ram[17062]  = 1;
  ram[17063]  = 1;
  ram[17064]  = 1;
  ram[17065]  = 1;
  ram[17066]  = 1;
  ram[17067]  = 1;
  ram[17068]  = 1;
  ram[17069]  = 1;
  ram[17070]  = 1;
  ram[17071]  = 1;
  ram[17072]  = 1;
  ram[17073]  = 1;
  ram[17074]  = 1;
  ram[17075]  = 1;
  ram[17076]  = 1;
  ram[17077]  = 1;
  ram[17078]  = 1;
  ram[17079]  = 1;
  ram[17080]  = 1;
  ram[17081]  = 1;
  ram[17082]  = 1;
  ram[17083]  = 1;
  ram[17084]  = 1;
  ram[17085]  = 1;
  ram[17086]  = 1;
  ram[17087]  = 1;
  ram[17088]  = 1;
  ram[17089]  = 1;
  ram[17090]  = 1;
  ram[17091]  = 1;
  ram[17092]  = 1;
  ram[17093]  = 1;
  ram[17094]  = 1;
  ram[17095]  = 1;
  ram[17096]  = 1;
  ram[17097]  = 1;
  ram[17098]  = 1;
  ram[17099]  = 1;
  ram[17100]  = 1;
  ram[17101]  = 1;
  ram[17102]  = 1;
  ram[17103]  = 1;
  ram[17104]  = 1;
  ram[17105]  = 1;
  ram[17106]  = 1;
  ram[17107]  = 1;
  ram[17108]  = 1;
  ram[17109]  = 1;
  ram[17110]  = 1;
  ram[17111]  = 1;
  ram[17112]  = 1;
  ram[17113]  = 1;
  ram[17114]  = 1;
  ram[17115]  = 1;
  ram[17116]  = 1;
  ram[17117]  = 1;
  ram[17118]  = 1;
  ram[17119]  = 1;
  ram[17120]  = 1;
  ram[17121]  = 1;
  ram[17122]  = 1;
  ram[17123]  = 1;
  ram[17124]  = 1;
  ram[17125]  = 1;
  ram[17126]  = 1;
  ram[17127]  = 1;
  ram[17128]  = 1;
  ram[17129]  = 1;
  ram[17130]  = 1;
  ram[17131]  = 1;
  ram[17132]  = 1;
  ram[17133]  = 1;
  ram[17134]  = 1;
  ram[17135]  = 1;
  ram[17136]  = 1;
  ram[17137]  = 1;
  ram[17138]  = 1;
  ram[17139]  = 1;
  ram[17140]  = 1;
  ram[17141]  = 1;
  ram[17142]  = 1;
  ram[17143]  = 1;
  ram[17144]  = 1;
  ram[17145]  = 1;
  ram[17146]  = 1;
  ram[17147]  = 1;
  ram[17148]  = 1;
  ram[17149]  = 1;
  ram[17150]  = 1;
  ram[17151]  = 1;
  ram[17152]  = 1;
  ram[17153]  = 1;
  ram[17154]  = 1;
  ram[17155]  = 1;
  ram[17156]  = 1;
  ram[17157]  = 1;
  ram[17158]  = 1;
  ram[17159]  = 1;
  ram[17160]  = 1;
  ram[17161]  = 1;
  ram[17162]  = 1;
  ram[17163]  = 1;
  ram[17164]  = 1;
  ram[17165]  = 1;
  ram[17166]  = 1;
  ram[17167]  = 1;
  ram[17168]  = 1;
  ram[17169]  = 1;
  ram[17170]  = 1;
  ram[17171]  = 1;
  ram[17172]  = 1;
  ram[17173]  = 1;
  ram[17174]  = 1;
  ram[17175]  = 1;
  ram[17176]  = 1;
  ram[17177]  = 1;
  ram[17178]  = 1;
  ram[17179]  = 1;
  ram[17180]  = 1;
  ram[17181]  = 1;
  ram[17182]  = 1;
  ram[17183]  = 1;
  ram[17184]  = 1;
  ram[17185]  = 1;
  ram[17186]  = 1;
  ram[17187]  = 1;
  ram[17188]  = 1;
  ram[17189]  = 1;
  ram[17190]  = 1;
  ram[17191]  = 1;
  ram[17192]  = 1;
  ram[17193]  = 1;
  ram[17194]  = 1;
  ram[17195]  = 1;
  ram[17196]  = 1;
  ram[17197]  = 1;
  ram[17198]  = 1;
  ram[17199]  = 1;
  ram[17200]  = 1;
  ram[17201]  = 1;
  ram[17202]  = 1;
  ram[17203]  = 1;
  ram[17204]  = 1;
  ram[17205]  = 1;
  ram[17206]  = 1;
  ram[17207]  = 1;
  ram[17208]  = 1;
  ram[17209]  = 1;
  ram[17210]  = 1;
  ram[17211]  = 1;
  ram[17212]  = 1;
  ram[17213]  = 1;
  ram[17214]  = 1;
  ram[17215]  = 1;
  ram[17216]  = 1;
  ram[17217]  = 1;
  ram[17218]  = 1;
  ram[17219]  = 1;
  ram[17220]  = 1;
  ram[17221]  = 1;
  ram[17222]  = 1;
  ram[17223]  = 1;
  ram[17224]  = 1;
  ram[17225]  = 1;
  ram[17226]  = 1;
  ram[17227]  = 1;
  ram[17228]  = 1;
  ram[17229]  = 1;
  ram[17230]  = 1;
  ram[17231]  = 1;
  ram[17232]  = 1;
  ram[17233]  = 1;
  ram[17234]  = 1;
  ram[17235]  = 1;
  ram[17236]  = 1;
  ram[17237]  = 1;
  ram[17238]  = 1;
  ram[17239]  = 1;
  ram[17240]  = 1;
  ram[17241]  = 1;
  ram[17242]  = 1;
  ram[17243]  = 1;
  ram[17244]  = 1;
  ram[17245]  = 1;
  ram[17246]  = 1;
  ram[17247]  = 1;
  ram[17248]  = 1;
  ram[17249]  = 1;
  ram[17250]  = 1;
  ram[17251]  = 1;
  ram[17252]  = 1;
  ram[17253]  = 1;
  ram[17254]  = 1;
  ram[17255]  = 1;
  ram[17256]  = 1;
  ram[17257]  = 1;
  ram[17258]  = 1;
  ram[17259]  = 1;
  ram[17260]  = 1;
  ram[17261]  = 1;
  ram[17262]  = 1;
  ram[17263]  = 1;
  ram[17264]  = 1;
  ram[17265]  = 1;
  ram[17266]  = 1;
  ram[17267]  = 1;
  ram[17268]  = 1;
  ram[17269]  = 1;
  ram[17270]  = 1;
  ram[17271]  = 1;
  ram[17272]  = 1;
  ram[17273]  = 1;
  ram[17274]  = 1;
  ram[17275]  = 1;
  ram[17276]  = 1;
  ram[17277]  = 1;
  ram[17278]  = 1;
  ram[17279]  = 1;
  ram[17280]  = 1;
  ram[17281]  = 1;
  ram[17282]  = 1;
  ram[17283]  = 1;
  ram[17284]  = 1;
  ram[17285]  = 1;
  ram[17286]  = 1;
  ram[17287]  = 1;
  ram[17288]  = 1;
  ram[17289]  = 1;
  ram[17290]  = 1;
  ram[17291]  = 1;
  ram[17292]  = 1;
  ram[17293]  = 1;
  ram[17294]  = 1;
  ram[17295]  = 1;
  ram[17296]  = 1;
  ram[17297]  = 1;
  ram[17298]  = 1;
  ram[17299]  = 1;
  ram[17300]  = 1;
  ram[17301]  = 1;
  ram[17302]  = 1;
  ram[17303]  = 1;
  ram[17304]  = 1;
  ram[17305]  = 1;
  ram[17306]  = 1;
  ram[17307]  = 1;
  ram[17308]  = 1;
  ram[17309]  = 1;
  ram[17310]  = 1;
  ram[17311]  = 1;
  ram[17312]  = 1;
  ram[17313]  = 1;
  ram[17314]  = 1;
  ram[17315]  = 1;
  ram[17316]  = 1;
  ram[17317]  = 1;
  ram[17318]  = 1;
  ram[17319]  = 1;
  ram[17320]  = 1;
  ram[17321]  = 1;
  ram[17322]  = 1;
  ram[17323]  = 1;
  ram[17324]  = 1;
  ram[17325]  = 1;
  ram[17326]  = 1;
  ram[17327]  = 1;
  ram[17328]  = 1;
  ram[17329]  = 1;
  ram[17330]  = 1;
  ram[17331]  = 1;
  ram[17332]  = 1;
  ram[17333]  = 1;
  ram[17334]  = 1;
  ram[17335]  = 1;
  ram[17336]  = 1;
  ram[17337]  = 1;
  ram[17338]  = 1;
  ram[17339]  = 1;
  ram[17340]  = 1;
  ram[17341]  = 1;
  ram[17342]  = 1;
  ram[17343]  = 1;
  ram[17344]  = 1;
  ram[17345]  = 1;
  ram[17346]  = 1;
  ram[17347]  = 1;
  ram[17348]  = 1;
  ram[17349]  = 1;
  ram[17350]  = 1;
  ram[17351]  = 1;
  ram[17352]  = 1;
  ram[17353]  = 1;
  ram[17354]  = 1;
  ram[17355]  = 1;
  ram[17356]  = 1;
  ram[17357]  = 1;
  ram[17358]  = 1;
  ram[17359]  = 1;
  ram[17360]  = 1;
  ram[17361]  = 1;
  ram[17362]  = 1;
  ram[17363]  = 1;
  ram[17364]  = 1;
  ram[17365]  = 1;
  ram[17366]  = 1;
  ram[17367]  = 1;
  ram[17368]  = 1;
  ram[17369]  = 1;
  ram[17370]  = 1;
  ram[17371]  = 1;
  ram[17372]  = 1;
  ram[17373]  = 1;
  ram[17374]  = 1;
  ram[17375]  = 1;
  ram[17376]  = 1;
  ram[17377]  = 1;
  ram[17378]  = 1;
  ram[17379]  = 1;
  ram[17380]  = 1;
  ram[17381]  = 1;
  ram[17382]  = 1;
  ram[17383]  = 1;
  ram[17384]  = 1;
  ram[17385]  = 1;
  ram[17386]  = 1;
  ram[17387]  = 1;
  ram[17388]  = 1;
  ram[17389]  = 1;
  ram[17390]  = 1;
  ram[17391]  = 1;
  ram[17392]  = 1;
  ram[17393]  = 1;
  ram[17394]  = 1;
  ram[17395]  = 1;
  ram[17396]  = 1;
  ram[17397]  = 1;
  ram[17398]  = 1;
  ram[17399]  = 1;
  ram[17400]  = 1;
  ram[17401]  = 1;
  ram[17402]  = 1;
  ram[17403]  = 1;
  ram[17404]  = 1;
  ram[17405]  = 1;
  ram[17406]  = 1;
  ram[17407]  = 1;
  ram[17408]  = 1;
  ram[17409]  = 1;
  ram[17410]  = 1;
  ram[17411]  = 1;
  ram[17412]  = 1;
  ram[17413]  = 1;
  ram[17414]  = 1;
  ram[17415]  = 1;
  ram[17416]  = 1;
  ram[17417]  = 1;
  ram[17418]  = 1;
  ram[17419]  = 1;
  ram[17420]  = 1;
  ram[17421]  = 1;
  ram[17422]  = 1;
  ram[17423]  = 1;
  ram[17424]  = 1;
  ram[17425]  = 1;
  ram[17426]  = 1;
  ram[17427]  = 1;
  ram[17428]  = 1;
  ram[17429]  = 1;
  ram[17430]  = 1;
  ram[17431]  = 1;
  ram[17432]  = 1;
  ram[17433]  = 1;
  ram[17434]  = 1;
  ram[17435]  = 1;
  ram[17436]  = 1;
  ram[17437]  = 1;
  ram[17438]  = 1;
  ram[17439]  = 1;
  ram[17440]  = 1;
  ram[17441]  = 1;
  ram[17442]  = 1;
  ram[17443]  = 1;
  ram[17444]  = 1;
  ram[17445]  = 1;
  ram[17446]  = 1;
  ram[17447]  = 1;
  ram[17448]  = 1;
  ram[17449]  = 1;
  ram[17450]  = 1;
  ram[17451]  = 1;
  ram[17452]  = 1;
  ram[17453]  = 1;
  ram[17454]  = 1;
  ram[17455]  = 1;
  ram[17456]  = 1;
  ram[17457]  = 1;
  ram[17458]  = 1;
  ram[17459]  = 1;
  ram[17460]  = 1;
  ram[17461]  = 1;
  ram[17462]  = 1;
  ram[17463]  = 1;
  ram[17464]  = 1;
  ram[17465]  = 1;
  ram[17466]  = 1;
  ram[17467]  = 1;
  ram[17468]  = 1;
  ram[17469]  = 1;
  ram[17470]  = 1;
  ram[17471]  = 1;
  ram[17472]  = 1;
  ram[17473]  = 1;
  ram[17474]  = 1;
  ram[17475]  = 1;
  ram[17476]  = 1;
  ram[17477]  = 1;
  ram[17478]  = 1;
  ram[17479]  = 1;
  ram[17480]  = 1;
  ram[17481]  = 1;
  ram[17482]  = 1;
  ram[17483]  = 1;
  ram[17484]  = 1;
  ram[17485]  = 1;
  ram[17486]  = 1;
  ram[17487]  = 1;
  ram[17488]  = 1;
  ram[17489]  = 1;
  ram[17490]  = 1;
  ram[17491]  = 1;
  ram[17492]  = 1;
  ram[17493]  = 1;
  ram[17494]  = 1;
  ram[17495]  = 1;
  ram[17496]  = 1;
  ram[17497]  = 1;
  ram[17498]  = 1;
  ram[17499]  = 1;
  ram[17500]  = 1;
  ram[17501]  = 1;
  ram[17502]  = 1;
  ram[17503]  = 1;
  ram[17504]  = 1;
  ram[17505]  = 1;
  ram[17506]  = 1;
  ram[17507]  = 1;
  ram[17508]  = 1;
  ram[17509]  = 1;
  ram[17510]  = 1;
  ram[17511]  = 1;
  ram[17512]  = 1;
  ram[17513]  = 1;
  ram[17514]  = 1;
  ram[17515]  = 1;
  ram[17516]  = 1;
  ram[17517]  = 1;
  ram[17518]  = 1;
  ram[17519]  = 1;
  ram[17520]  = 1;
  ram[17521]  = 1;
  ram[17522]  = 1;
  ram[17523]  = 1;
  ram[17524]  = 1;
  ram[17525]  = 1;
  ram[17526]  = 1;
  ram[17527]  = 1;
  ram[17528]  = 1;
  ram[17529]  = 1;
  ram[17530]  = 1;
  ram[17531]  = 1;
  ram[17532]  = 1;
  ram[17533]  = 1;
  ram[17534]  = 1;
  ram[17535]  = 1;
  ram[17536]  = 1;
  ram[17537]  = 1;
  ram[17538]  = 1;
  ram[17539]  = 1;
  ram[17540]  = 1;
  ram[17541]  = 1;
  ram[17542]  = 1;
  ram[17543]  = 1;
  ram[17544]  = 1;
  ram[17545]  = 1;
  ram[17546]  = 1;
  ram[17547]  = 1;
  ram[17548]  = 1;
  ram[17549]  = 1;
  ram[17550]  = 1;
  ram[17551]  = 1;
  ram[17552]  = 1;
  ram[17553]  = 1;
  ram[17554]  = 1;
  ram[17555]  = 1;
  ram[17556]  = 1;
  ram[17557]  = 1;
  ram[17558]  = 1;
  ram[17559]  = 1;
  ram[17560]  = 1;
  ram[17561]  = 1;
  ram[17562]  = 1;
  ram[17563]  = 1;
  ram[17564]  = 1;
  ram[17565]  = 1;
  ram[17566]  = 1;
  ram[17567]  = 1;
  ram[17568]  = 1;
  ram[17569]  = 1;
  ram[17570]  = 1;
  ram[17571]  = 1;
  ram[17572]  = 1;
  ram[17573]  = 1;
  ram[17574]  = 1;
  ram[17575]  = 1;
  ram[17576]  = 1;
  ram[17577]  = 1;
  ram[17578]  = 1;
  ram[17579]  = 1;
  ram[17580]  = 1;
  ram[17581]  = 1;
  ram[17582]  = 1;
  ram[17583]  = 1;
  ram[17584]  = 1;
  ram[17585]  = 1;
  ram[17586]  = 1;
  ram[17587]  = 1;
  ram[17588]  = 1;
  ram[17589]  = 1;
  ram[17590]  = 1;
  ram[17591]  = 1;
  ram[17592]  = 1;
  ram[17593]  = 1;
  ram[17594]  = 1;
  ram[17595]  = 1;
  ram[17596]  = 1;
  ram[17597]  = 1;
  ram[17598]  = 1;
  ram[17599]  = 1;
  ram[17600]  = 1;
  ram[17601]  = 1;
  ram[17602]  = 1;
  ram[17603]  = 1;
  ram[17604]  = 1;
  ram[17605]  = 1;
  ram[17606]  = 1;
  ram[17607]  = 1;
  ram[17608]  = 1;
  ram[17609]  = 1;
  ram[17610]  = 1;
  ram[17611]  = 1;
  ram[17612]  = 1;
  ram[17613]  = 1;
  ram[17614]  = 1;
  ram[17615]  = 1;
  ram[17616]  = 1;
  ram[17617]  = 1;
  ram[17618]  = 1;
  ram[17619]  = 1;
  ram[17620]  = 1;
  ram[17621]  = 1;
  ram[17622]  = 1;
  ram[17623]  = 1;
  ram[17624]  = 1;
  ram[17625]  = 1;
  ram[17626]  = 1;
  ram[17627]  = 1;
  ram[17628]  = 1;
  ram[17629]  = 1;
  ram[17630]  = 1;
  ram[17631]  = 1;
  ram[17632]  = 1;
  ram[17633]  = 1;
  ram[17634]  = 1;
  ram[17635]  = 1;
  ram[17636]  = 1;
  ram[17637]  = 1;
  ram[17638]  = 1;
  ram[17639]  = 1;
  ram[17640]  = 1;
  ram[17641]  = 1;
  ram[17642]  = 1;
  ram[17643]  = 1;
  ram[17644]  = 1;
  ram[17645]  = 1;
  ram[17646]  = 1;
  ram[17647]  = 1;
  ram[17648]  = 1;
  ram[17649]  = 1;
  ram[17650]  = 1;
  ram[17651]  = 1;
  ram[17652]  = 1;
  ram[17653]  = 1;
  ram[17654]  = 1;
  ram[17655]  = 1;
  ram[17656]  = 1;
  ram[17657]  = 1;
  ram[17658]  = 1;
  ram[17659]  = 1;
  ram[17660]  = 1;
  ram[17661]  = 1;
  ram[17662]  = 1;
  ram[17663]  = 1;
  ram[17664]  = 1;
  ram[17665]  = 1;
  ram[17666]  = 1;
  ram[17667]  = 1;
  ram[17668]  = 1;
  ram[17669]  = 1;
  ram[17670]  = 1;
  ram[17671]  = 1;
  ram[17672]  = 1;
  ram[17673]  = 1;
  ram[17674]  = 1;
  ram[17675]  = 1;
  ram[17676]  = 1;
  ram[17677]  = 1;
  ram[17678]  = 1;
  ram[17679]  = 1;
  ram[17680]  = 1;
  ram[17681]  = 1;
  ram[17682]  = 1;
  ram[17683]  = 1;
  ram[17684]  = 1;
  ram[17685]  = 1;
  ram[17686]  = 1;
  ram[17687]  = 1;
  ram[17688]  = 1;
  ram[17689]  = 1;
  ram[17690]  = 1;
  ram[17691]  = 1;
  ram[17692]  = 1;
  ram[17693]  = 1;
  ram[17694]  = 1;
  ram[17695]  = 1;
  ram[17696]  = 1;
  ram[17697]  = 1;
  ram[17698]  = 1;
  ram[17699]  = 1;
  ram[17700]  = 1;
  ram[17701]  = 1;
  ram[17702]  = 1;
  ram[17703]  = 1;
  ram[17704]  = 1;
  ram[17705]  = 1;
  ram[17706]  = 1;
  ram[17707]  = 1;
  ram[17708]  = 1;
  ram[17709]  = 1;
  ram[17710]  = 1;
  ram[17711]  = 1;
  ram[17712]  = 1;
  ram[17713]  = 1;
  ram[17714]  = 1;
  ram[17715]  = 1;
  ram[17716]  = 1;
  ram[17717]  = 1;
  ram[17718]  = 1;
  ram[17719]  = 1;
  ram[17720]  = 1;
  ram[17721]  = 1;
  ram[17722]  = 1;
  ram[17723]  = 1;
  ram[17724]  = 1;
  ram[17725]  = 1;
  ram[17726]  = 1;
  ram[17727]  = 1;
  ram[17728]  = 1;
  ram[17729]  = 1;
  ram[17730]  = 1;
  ram[17731]  = 1;
  ram[17732]  = 1;
  ram[17733]  = 1;
  ram[17734]  = 1;
  ram[17735]  = 1;
  ram[17736]  = 1;
  ram[17737]  = 1;
  ram[17738]  = 1;
  ram[17739]  = 1;
  ram[17740]  = 1;
  ram[17741]  = 1;
  ram[17742]  = 1;
  ram[17743]  = 1;
  ram[17744]  = 1;
  ram[17745]  = 1;
  ram[17746]  = 1;
  ram[17747]  = 1;
  ram[17748]  = 1;
  ram[17749]  = 1;
  ram[17750]  = 1;
  ram[17751]  = 1;
  ram[17752]  = 1;
  ram[17753]  = 1;
  ram[17754]  = 1;
  ram[17755]  = 1;
  ram[17756]  = 1;
  ram[17757]  = 1;
  ram[17758]  = 1;
  ram[17759]  = 1;
  ram[17760]  = 1;
  ram[17761]  = 1;
  ram[17762]  = 1;
  ram[17763]  = 1;
  ram[17764]  = 1;
  ram[17765]  = 1;
  ram[17766]  = 1;
  ram[17767]  = 1;
  ram[17768]  = 1;
  ram[17769]  = 1;
  ram[17770]  = 1;
  ram[17771]  = 1;
  ram[17772]  = 1;
  ram[17773]  = 1;
  ram[17774]  = 1;
  ram[17775]  = 1;
  ram[17776]  = 1;
  ram[17777]  = 1;
  ram[17778]  = 1;
  ram[17779]  = 1;
  ram[17780]  = 1;
  ram[17781]  = 1;
  ram[17782]  = 1;
  ram[17783]  = 1;
  ram[17784]  = 1;
  ram[17785]  = 1;
  ram[17786]  = 1;
  ram[17787]  = 1;
  ram[17788]  = 1;
  ram[17789]  = 1;
  ram[17790]  = 1;
  ram[17791]  = 1;
  ram[17792]  = 1;
  ram[17793]  = 1;
  ram[17794]  = 1;
  ram[17795]  = 1;
  ram[17796]  = 1;
  ram[17797]  = 1;
  ram[17798]  = 1;
  ram[17799]  = 1;
  ram[17800]  = 1;
  ram[17801]  = 1;
  ram[17802]  = 1;
  ram[17803]  = 1;
  ram[17804]  = 1;
  ram[17805]  = 1;
  ram[17806]  = 1;
  ram[17807]  = 1;
  ram[17808]  = 1;
  ram[17809]  = 1;
  ram[17810]  = 1;
  ram[17811]  = 1;
  ram[17812]  = 1;
  ram[17813]  = 1;
  ram[17814]  = 1;
  ram[17815]  = 1;
  ram[17816]  = 1;
  ram[17817]  = 1;
  ram[17818]  = 1;
  ram[17819]  = 1;
  ram[17820]  = 1;
  ram[17821]  = 1;
  ram[17822]  = 1;
  ram[17823]  = 1;
  ram[17824]  = 1;
  ram[17825]  = 1;
  ram[17826]  = 1;
  ram[17827]  = 1;
  ram[17828]  = 1;
  ram[17829]  = 1;
  ram[17830]  = 1;
  ram[17831]  = 1;
  ram[17832]  = 1;
  ram[17833]  = 1;
  ram[17834]  = 1;
  ram[17835]  = 1;
  ram[17836]  = 1;
  ram[17837]  = 1;
  ram[17838]  = 1;
  ram[17839]  = 1;
  ram[17840]  = 1;
  ram[17841]  = 1;
  ram[17842]  = 1;
  ram[17843]  = 1;
  ram[17844]  = 1;
  ram[17845]  = 1;
  ram[17846]  = 1;
  ram[17847]  = 1;
  ram[17848]  = 1;
  ram[17849]  = 1;
  ram[17850]  = 1;
  ram[17851]  = 1;
  ram[17852]  = 1;
  ram[17853]  = 1;
  ram[17854]  = 1;
  ram[17855]  = 1;
  ram[17856]  = 1;
  ram[17857]  = 1;
  ram[17858]  = 1;
  ram[17859]  = 1;
  ram[17860]  = 1;
  ram[17861]  = 1;
  ram[17862]  = 1;
  ram[17863]  = 1;
  ram[17864]  = 1;
  ram[17865]  = 1;
  ram[17866]  = 1;
  ram[17867]  = 1;
  ram[17868]  = 1;
  ram[17869]  = 1;
  ram[17870]  = 1;
  ram[17871]  = 1;
  ram[17872]  = 1;
  ram[17873]  = 1;
  ram[17874]  = 1;
  ram[17875]  = 1;
  ram[17876]  = 1;
  ram[17877]  = 1;
  ram[17878]  = 1;
  ram[17879]  = 1;
  ram[17880]  = 1;
  ram[17881]  = 1;
  ram[17882]  = 1;
  ram[17883]  = 1;
  ram[17884]  = 1;
  ram[17885]  = 1;
  ram[17886]  = 1;
  ram[17887]  = 1;
  ram[17888]  = 1;
  ram[17889]  = 1;
  ram[17890]  = 1;
  ram[17891]  = 1;
  ram[17892]  = 1;
  ram[17893]  = 1;
  ram[17894]  = 1;
  ram[17895]  = 1;
  ram[17896]  = 1;
  ram[17897]  = 1;
  ram[17898]  = 1;
  ram[17899]  = 1;
  ram[17900]  = 1;
  ram[17901]  = 1;
  ram[17902]  = 1;
  ram[17903]  = 1;
  ram[17904]  = 1;
  ram[17905]  = 1;
  ram[17906]  = 1;
  ram[17907]  = 1;
  ram[17908]  = 1;
  ram[17909]  = 1;
  ram[17910]  = 1;
  ram[17911]  = 1;
  ram[17912]  = 1;
  ram[17913]  = 1;
  ram[17914]  = 1;
  ram[17915]  = 1;
  ram[17916]  = 1;
  ram[17917]  = 1;
  ram[17918]  = 1;
  ram[17919]  = 1;
  ram[17920]  = 1;
  ram[17921]  = 1;
  ram[17922]  = 1;
  ram[17923]  = 1;
  ram[17924]  = 1;
  ram[17925]  = 1;
  ram[17926]  = 1;
  ram[17927]  = 1;
  ram[17928]  = 1;
  ram[17929]  = 1;
  ram[17930]  = 1;
  ram[17931]  = 1;
  ram[17932]  = 1;
  ram[17933]  = 1;
  ram[17934]  = 1;
  ram[17935]  = 1;
  ram[17936]  = 1;
  ram[17937]  = 1;
  ram[17938]  = 1;
  ram[17939]  = 1;
  ram[17940]  = 1;
  ram[17941]  = 1;
  ram[17942]  = 1;
  ram[17943]  = 1;
  ram[17944]  = 1;
  ram[17945]  = 1;
  ram[17946]  = 1;
  ram[17947]  = 1;
  ram[17948]  = 1;
  ram[17949]  = 1;
  ram[17950]  = 1;
  ram[17951]  = 1;
  ram[17952]  = 1;
  ram[17953]  = 1;
  ram[17954]  = 1;
  ram[17955]  = 1;
  ram[17956]  = 1;
  ram[17957]  = 1;
  ram[17958]  = 1;
  ram[17959]  = 1;
  ram[17960]  = 1;
  ram[17961]  = 1;
  ram[17962]  = 1;
  ram[17963]  = 1;
  ram[17964]  = 1;
  ram[17965]  = 1;
  ram[17966]  = 1;
  ram[17967]  = 1;
  ram[17968]  = 1;
  ram[17969]  = 1;
  ram[17970]  = 1;
  ram[17971]  = 1;
  ram[17972]  = 1;
  ram[17973]  = 1;
  ram[17974]  = 1;
  ram[17975]  = 1;
  ram[17976]  = 1;
  ram[17977]  = 1;
  ram[17978]  = 1;
  ram[17979]  = 1;
  ram[17980]  = 1;
  ram[17981]  = 1;
  ram[17982]  = 1;
  ram[17983]  = 1;
  ram[17984]  = 1;
  ram[17985]  = 1;
  ram[17986]  = 1;
  ram[17987]  = 1;
  ram[17988]  = 1;
  ram[17989]  = 1;
  ram[17990]  = 1;
  ram[17991]  = 1;
  ram[17992]  = 1;
  ram[17993]  = 1;
  ram[17994]  = 1;
  ram[17995]  = 1;
  ram[17996]  = 1;
  ram[17997]  = 1;
  ram[17998]  = 1;
  ram[17999]  = 1;
  ram[18000]  = 1;
  ram[18001]  = 1;
  ram[18002]  = 1;
  ram[18003]  = 1;
  ram[18004]  = 1;
  ram[18005]  = 1;
  ram[18006]  = 1;
  ram[18007]  = 1;
  ram[18008]  = 1;
  ram[18009]  = 1;
  ram[18010]  = 1;
  ram[18011]  = 1;
  ram[18012]  = 1;
  ram[18013]  = 1;
  ram[18014]  = 1;
  ram[18015]  = 1;
  ram[18016]  = 1;
  ram[18017]  = 1;
  ram[18018]  = 1;
  ram[18019]  = 1;
  ram[18020]  = 1;
  ram[18021]  = 1;
  ram[18022]  = 1;
  ram[18023]  = 1;
  ram[18024]  = 1;
  ram[18025]  = 1;
  ram[18026]  = 1;
  ram[18027]  = 1;
  ram[18028]  = 1;
  ram[18029]  = 1;
  ram[18030]  = 1;
  ram[18031]  = 1;
  ram[18032]  = 1;
  ram[18033]  = 1;
  ram[18034]  = 1;
  ram[18035]  = 1;
  ram[18036]  = 1;
  ram[18037]  = 1;
  ram[18038]  = 1;
  ram[18039]  = 1;
  ram[18040]  = 1;
  ram[18041]  = 1;
  ram[18042]  = 1;
  ram[18043]  = 1;
  ram[18044]  = 1;
  ram[18045]  = 1;
  ram[18046]  = 1;
  ram[18047]  = 1;
  ram[18048]  = 1;
  ram[18049]  = 1;
  ram[18050]  = 1;
  ram[18051]  = 1;
  ram[18052]  = 1;
  ram[18053]  = 1;
  ram[18054]  = 1;
  ram[18055]  = 1;
  ram[18056]  = 1;
  ram[18057]  = 1;
  ram[18058]  = 1;
  ram[18059]  = 1;
  ram[18060]  = 1;
  ram[18061]  = 1;
  ram[18062]  = 1;
  ram[18063]  = 1;
  ram[18064]  = 1;
  ram[18065]  = 1;
  ram[18066]  = 1;
  ram[18067]  = 1;
  ram[18068]  = 1;
  ram[18069]  = 1;
  ram[18070]  = 1;
  ram[18071]  = 1;
  ram[18072]  = 1;
  ram[18073]  = 1;
  ram[18074]  = 1;
  ram[18075]  = 1;
  ram[18076]  = 1;
  ram[18077]  = 1;
  ram[18078]  = 1;
  ram[18079]  = 1;
  ram[18080]  = 1;
  ram[18081]  = 1;
  ram[18082]  = 1;
  ram[18083]  = 1;
  ram[18084]  = 1;
  ram[18085]  = 1;
  ram[18086]  = 1;
  ram[18087]  = 1;
  ram[18088]  = 1;
  ram[18089]  = 1;
  ram[18090]  = 1;
  ram[18091]  = 1;
  ram[18092]  = 1;
  ram[18093]  = 1;
  ram[18094]  = 1;
  ram[18095]  = 1;
  ram[18096]  = 1;
  ram[18097]  = 0;
  ram[18098]  = 1;
  ram[18099]  = 1;
  ram[18100]  = 1;
  ram[18101]  = 1;
  ram[18102]  = 1;
  ram[18103]  = 1;
  ram[18104]  = 1;
  ram[18105]  = 1;
  ram[18106]  = 1;
  ram[18107]  = 1;
  ram[18108]  = 1;
  ram[18109]  = 1;
  ram[18110]  = 1;
  ram[18111]  = 1;
  ram[18112]  = 1;
  ram[18113]  = 1;
  ram[18114]  = 1;
  ram[18115]  = 1;
  ram[18116]  = 1;
  ram[18117]  = 1;
  ram[18118]  = 1;
  ram[18119]  = 1;
  ram[18120]  = 1;
  ram[18121]  = 1;
  ram[18122]  = 1;
  ram[18123]  = 1;
  ram[18124]  = 1;
  ram[18125]  = 1;
  ram[18126]  = 1;
  ram[18127]  = 1;
  ram[18128]  = 1;
  ram[18129]  = 1;
  ram[18130]  = 1;
  ram[18131]  = 1;
  ram[18132]  = 1;
  ram[18133]  = 1;
  ram[18134]  = 1;
  ram[18135]  = 1;
  ram[18136]  = 1;
  ram[18137]  = 1;
  ram[18138]  = 1;
  ram[18139]  = 1;
  ram[18140]  = 1;
  ram[18141]  = 1;
  ram[18142]  = 1;
  ram[18143]  = 1;
  ram[18144]  = 1;
  ram[18145]  = 1;
  ram[18146]  = 1;
  ram[18147]  = 1;
  ram[18148]  = 1;
  ram[18149]  = 1;
  ram[18150]  = 1;
  ram[18151]  = 1;
  ram[18152]  = 1;
  ram[18153]  = 1;
  ram[18154]  = 1;
  ram[18155]  = 1;
  ram[18156]  = 1;
  ram[18157]  = 1;
  ram[18158]  = 1;
  ram[18159]  = 1;
  ram[18160]  = 1;
  ram[18161]  = 1;
  ram[18162]  = 1;
  ram[18163]  = 1;
  ram[18164]  = 1;
  ram[18165]  = 1;
  ram[18166]  = 1;
  ram[18167]  = 1;
  ram[18168]  = 1;
  ram[18169]  = 1;
  ram[18170]  = 1;
  ram[18171]  = 1;
  ram[18172]  = 1;
  ram[18173]  = 1;
  ram[18174]  = 1;
  ram[18175]  = 1;
  ram[18176]  = 1;
  ram[18177]  = 1;
  ram[18178]  = 1;
  ram[18179]  = 1;
  ram[18180]  = 1;
  ram[18181]  = 1;
  ram[18182]  = 1;
  ram[18183]  = 1;
  ram[18184]  = 1;
  ram[18185]  = 1;
  ram[18186]  = 1;
  ram[18187]  = 1;
  ram[18188]  = 1;
  ram[18189]  = 1;
  ram[18190]  = 1;
  ram[18191]  = 1;
  ram[18192]  = 1;
  ram[18193]  = 1;
  ram[18194]  = 1;
  ram[18195]  = 1;
  ram[18196]  = 1;
  ram[18197]  = 1;
  ram[18198]  = 1;
  ram[18199]  = 1;
  ram[18200]  = 1;
  ram[18201]  = 1;
  ram[18202]  = 1;
  ram[18203]  = 1;
  ram[18204]  = 1;
  ram[18205]  = 1;
  ram[18206]  = 1;
  ram[18207]  = 1;
  ram[18208]  = 1;
  ram[18209]  = 1;
  ram[18210]  = 1;
  ram[18211]  = 1;
  ram[18212]  = 1;
  ram[18213]  = 1;
  ram[18214]  = 1;
  ram[18215]  = 1;
  ram[18216]  = 1;
  ram[18217]  = 1;
  ram[18218]  = 1;
  ram[18219]  = 1;
  ram[18220]  = 1;
  ram[18221]  = 1;
  ram[18222]  = 1;
  ram[18223]  = 1;
  ram[18224]  = 1;
  ram[18225]  = 1;
  ram[18226]  = 1;
  ram[18227]  = 1;
  ram[18228]  = 1;
  ram[18229]  = 1;
  ram[18230]  = 1;
  ram[18231]  = 1;
  ram[18232]  = 1;
  ram[18233]  = 1;
  ram[18234]  = 1;
  ram[18235]  = 1;
  ram[18236]  = 1;
  ram[18237]  = 1;
  ram[18238]  = 1;
  ram[18239]  = 1;
  ram[18240]  = 1;
  ram[18241]  = 1;
  ram[18242]  = 1;
  ram[18243]  = 1;
  ram[18244]  = 1;
  ram[18245]  = 1;
  ram[18246]  = 1;
  ram[18247]  = 1;
  ram[18248]  = 1;
  ram[18249]  = 1;
  ram[18250]  = 1;
  ram[18251]  = 1;
  ram[18252]  = 1;
  ram[18253]  = 1;
  ram[18254]  = 1;
  ram[18255]  = 1;
  ram[18256]  = 1;
  ram[18257]  = 1;
  ram[18258]  = 1;
  ram[18259]  = 1;
  ram[18260]  = 1;
  ram[18261]  = 1;
  ram[18262]  = 1;
  ram[18263]  = 1;
  ram[18264]  = 1;
  ram[18265]  = 1;
  ram[18266]  = 1;
  ram[18267]  = 1;
  ram[18268]  = 1;
  ram[18269]  = 1;
  ram[18270]  = 1;
  ram[18271]  = 1;
  ram[18272]  = 1;
  ram[18273]  = 1;
  ram[18274]  = 1;
  ram[18275]  = 1;
  ram[18276]  = 1;
  ram[18277]  = 1;
  ram[18278]  = 1;
  ram[18279]  = 1;
  ram[18280]  = 1;
  ram[18281]  = 1;
  ram[18282]  = 1;
  ram[18283]  = 1;
  ram[18284]  = 1;
  ram[18285]  = 1;
  ram[18286]  = 1;
  ram[18287]  = 1;
  ram[18288]  = 1;
  ram[18289]  = 1;
  ram[18290]  = 1;
  ram[18291]  = 1;
  ram[18292]  = 1;
  ram[18293]  = 1;
  ram[18294]  = 1;
  ram[18295]  = 1;
  ram[18296]  = 1;
  ram[18297]  = 1;
  ram[18298]  = 1;
  ram[18299]  = 1;
  ram[18300]  = 1;
  ram[18301]  = 1;
  ram[18302]  = 1;
  ram[18303]  = 1;
  ram[18304]  = 1;
  ram[18305]  = 1;
  ram[18306]  = 1;
  ram[18307]  = 1;
  ram[18308]  = 1;
  ram[18309]  = 1;
  ram[18310]  = 1;
  ram[18311]  = 1;
  ram[18312]  = 1;
  ram[18313]  = 1;
  ram[18314]  = 1;
  ram[18315]  = 1;
  ram[18316]  = 1;
  ram[18317]  = 1;
  ram[18318]  = 1;
  ram[18319]  = 1;
  ram[18320]  = 1;
  ram[18321]  = 1;
  ram[18322]  = 1;
  ram[18323]  = 1;
  ram[18324]  = 1;
  ram[18325]  = 1;
  ram[18326]  = 1;
  ram[18327]  = 1;
  ram[18328]  = 1;
  ram[18329]  = 1;
  ram[18330]  = 1;
  ram[18331]  = 1;
  ram[18332]  = 1;
  ram[18333]  = 1;
  ram[18334]  = 1;
  ram[18335]  = 1;
  ram[18336]  = 1;
  ram[18337]  = 1;
  ram[18338]  = 1;
  ram[18339]  = 1;
  ram[18340]  = 1;
  ram[18341]  = 1;
  ram[18342]  = 1;
  ram[18343]  = 1;
  ram[18344]  = 1;
  ram[18345]  = 0;
  ram[18346]  = 0;
  ram[18347]  = 0;
  ram[18348]  = 0;
  ram[18349]  = 0;
  ram[18350]  = 0;
  ram[18351]  = 1;
  ram[18352]  = 1;
  ram[18353]  = 1;
  ram[18354]  = 1;
  ram[18355]  = 1;
  ram[18356]  = 1;
  ram[18357]  = 1;
  ram[18358]  = 1;
  ram[18359]  = 1;
  ram[18360]  = 1;
  ram[18361]  = 1;
  ram[18362]  = 1;
  ram[18363]  = 1;
  ram[18364]  = 1;
  ram[18365]  = 1;
  ram[18366]  = 1;
  ram[18367]  = 1;
  ram[18368]  = 1;
  ram[18369]  = 1;
  ram[18370]  = 1;
  ram[18371]  = 1;
  ram[18372]  = 1;
  ram[18373]  = 1;
  ram[18374]  = 1;
  ram[18375]  = 1;
  ram[18376]  = 1;
  ram[18377]  = 1;
  ram[18378]  = 1;
  ram[18379]  = 1;
  ram[18380]  = 1;
  ram[18381]  = 1;
  ram[18382]  = 1;
  ram[18383]  = 1;
  ram[18384]  = 1;
  ram[18385]  = 1;
  ram[18386]  = 1;
  ram[18387]  = 1;
  ram[18388]  = 1;
  ram[18389]  = 1;
  ram[18390]  = 1;
  ram[18391]  = 1;
  ram[18392]  = 1;
  ram[18393]  = 1;
  ram[18394]  = 1;
  ram[18395]  = 1;
  ram[18396]  = 1;
  ram[18397]  = 0;
  ram[18398]  = 1;
  ram[18399]  = 1;
  ram[18400]  = 1;
  ram[18401]  = 1;
  ram[18402]  = 1;
  ram[18403]  = 1;
  ram[18404]  = 1;
  ram[18405]  = 1;
  ram[18406]  = 1;
  ram[18407]  = 1;
  ram[18408]  = 1;
  ram[18409]  = 1;
  ram[18410]  = 1;
  ram[18411]  = 1;
  ram[18412]  = 1;
  ram[18413]  = 1;
  ram[18414]  = 1;
  ram[18415]  = 1;
  ram[18416]  = 1;
  ram[18417]  = 1;
  ram[18418]  = 1;
  ram[18419]  = 1;
  ram[18420]  = 1;
  ram[18421]  = 1;
  ram[18422]  = 0;
  ram[18423]  = 0;
  ram[18424]  = 0;
  ram[18425]  = 0;
  ram[18426]  = 0;
  ram[18427]  = 1;
  ram[18428]  = 1;
  ram[18429]  = 1;
  ram[18430]  = 1;
  ram[18431]  = 1;
  ram[18432]  = 1;
  ram[18433]  = 1;
  ram[18434]  = 1;
  ram[18435]  = 1;
  ram[18436]  = 1;
  ram[18437]  = 1;
  ram[18438]  = 1;
  ram[18439]  = 1;
  ram[18440]  = 1;
  ram[18441]  = 1;
  ram[18442]  = 1;
  ram[18443]  = 1;
  ram[18444]  = 1;
  ram[18445]  = 1;
  ram[18446]  = 1;
  ram[18447]  = 1;
  ram[18448]  = 1;
  ram[18449]  = 1;
  ram[18450]  = 1;
  ram[18451]  = 1;
  ram[18452]  = 1;
  ram[18453]  = 1;
  ram[18454]  = 1;
  ram[18455]  = 1;
  ram[18456]  = 1;
  ram[18457]  = 1;
  ram[18458]  = 1;
  ram[18459]  = 1;
  ram[18460]  = 1;
  ram[18461]  = 1;
  ram[18462]  = 1;
  ram[18463]  = 1;
  ram[18464]  = 1;
  ram[18465]  = 1;
  ram[18466]  = 1;
  ram[18467]  = 1;
  ram[18468]  = 1;
  ram[18469]  = 1;
  ram[18470]  = 1;
  ram[18471]  = 1;
  ram[18472]  = 1;
  ram[18473]  = 1;
  ram[18474]  = 1;
  ram[18475]  = 1;
  ram[18476]  = 1;
  ram[18477]  = 1;
  ram[18478]  = 1;
  ram[18479]  = 1;
  ram[18480]  = 1;
  ram[18481]  = 1;
  ram[18482]  = 1;
  ram[18483]  = 1;
  ram[18484]  = 1;
  ram[18485]  = 1;
  ram[18486]  = 1;
  ram[18487]  = 1;
  ram[18488]  = 1;
  ram[18489]  = 1;
  ram[18490]  = 1;
  ram[18491]  = 1;
  ram[18492]  = 1;
  ram[18493]  = 1;
  ram[18494]  = 1;
  ram[18495]  = 1;
  ram[18496]  = 1;
  ram[18497]  = 1;
  ram[18498]  = 1;
  ram[18499]  = 1;
  ram[18500]  = 1;
  ram[18501]  = 1;
  ram[18502]  = 1;
  ram[18503]  = 1;
  ram[18504]  = 1;
  ram[18505]  = 1;
  ram[18506]  = 1;
  ram[18507]  = 1;
  ram[18508]  = 1;
  ram[18509]  = 1;
  ram[18510]  = 1;
  ram[18511]  = 1;
  ram[18512]  = 1;
  ram[18513]  = 1;
  ram[18514]  = 1;
  ram[18515]  = 1;
  ram[18516]  = 1;
  ram[18517]  = 1;
  ram[18518]  = 1;
  ram[18519]  = 1;
  ram[18520]  = 1;
  ram[18521]  = 1;
  ram[18522]  = 1;
  ram[18523]  = 1;
  ram[18524]  = 1;
  ram[18525]  = 1;
  ram[18526]  = 1;
  ram[18527]  = 1;
  ram[18528]  = 1;
  ram[18529]  = 1;
  ram[18530]  = 1;
  ram[18531]  = 1;
  ram[18532]  = 1;
  ram[18533]  = 1;
  ram[18534]  = 1;
  ram[18535]  = 1;
  ram[18536]  = 1;
  ram[18537]  = 1;
  ram[18538]  = 1;
  ram[18539]  = 1;
  ram[18540]  = 1;
  ram[18541]  = 1;
  ram[18542]  = 1;
  ram[18543]  = 1;
  ram[18544]  = 1;
  ram[18545]  = 1;
  ram[18546]  = 1;
  ram[18547]  = 1;
  ram[18548]  = 1;
  ram[18549]  = 1;
  ram[18550]  = 1;
  ram[18551]  = 1;
  ram[18552]  = 1;
  ram[18553]  = 1;
  ram[18554]  = 1;
  ram[18555]  = 1;
  ram[18556]  = 1;
  ram[18557]  = 1;
  ram[18558]  = 1;
  ram[18559]  = 1;
  ram[18560]  = 1;
  ram[18561]  = 1;
  ram[18562]  = 1;
  ram[18563]  = 1;
  ram[18564]  = 1;
  ram[18565]  = 1;
  ram[18566]  = 1;
  ram[18567]  = 1;
  ram[18568]  = 1;
  ram[18569]  = 1;
  ram[18570]  = 1;
  ram[18571]  = 1;
  ram[18572]  = 1;
  ram[18573]  = 1;
  ram[18574]  = 1;
  ram[18575]  = 1;
  ram[18576]  = 1;
  ram[18577]  = 1;
  ram[18578]  = 1;
  ram[18579]  = 1;
  ram[18580]  = 1;
  ram[18581]  = 1;
  ram[18582]  = 1;
  ram[18583]  = 1;
  ram[18584]  = 1;
  ram[18585]  = 1;
  ram[18586]  = 1;
  ram[18587]  = 1;
  ram[18588]  = 1;
  ram[18589]  = 1;
  ram[18590]  = 1;
  ram[18591]  = 1;
  ram[18592]  = 1;
  ram[18593]  = 1;
  ram[18594]  = 1;
  ram[18595]  = 1;
  ram[18596]  = 1;
  ram[18597]  = 1;
  ram[18598]  = 1;
  ram[18599]  = 1;
  ram[18600]  = 1;
  ram[18601]  = 1;
  ram[18602]  = 1;
  ram[18603]  = 1;
  ram[18604]  = 1;
  ram[18605]  = 1;
  ram[18606]  = 1;
  ram[18607]  = 1;
  ram[18608]  = 1;
  ram[18609]  = 1;
  ram[18610]  = 1;
  ram[18611]  = 1;
  ram[18612]  = 1;
  ram[18613]  = 1;
  ram[18614]  = 1;
  ram[18615]  = 1;
  ram[18616]  = 1;
  ram[18617]  = 1;
  ram[18618]  = 1;
  ram[18619]  = 1;
  ram[18620]  = 1;
  ram[18621]  = 1;
  ram[18622]  = 1;
  ram[18623]  = 1;
  ram[18624]  = 1;
  ram[18625]  = 1;
  ram[18626]  = 1;
  ram[18627]  = 1;
  ram[18628]  = 1;
  ram[18629]  = 1;
  ram[18630]  = 1;
  ram[18631]  = 1;
  ram[18632]  = 1;
  ram[18633]  = 1;
  ram[18634]  = 1;
  ram[18635]  = 1;
  ram[18636]  = 1;
  ram[18637]  = 1;
  ram[18638]  = 1;
  ram[18639]  = 1;
  ram[18640]  = 1;
  ram[18641]  = 1;
  ram[18642]  = 1;
  ram[18643]  = 1;
  ram[18644]  = 1;
  ram[18645]  = 0;
  ram[18646]  = 0;
  ram[18647]  = 0;
  ram[18648]  = 0;
  ram[18649]  = 0;
  ram[18650]  = 0;
  ram[18651]  = 1;
  ram[18652]  = 1;
  ram[18653]  = 1;
  ram[18654]  = 1;
  ram[18655]  = 1;
  ram[18656]  = 1;
  ram[18657]  = 1;
  ram[18658]  = 1;
  ram[18659]  = 1;
  ram[18660]  = 1;
  ram[18661]  = 1;
  ram[18662]  = 1;
  ram[18663]  = 1;
  ram[18664]  = 1;
  ram[18665]  = 1;
  ram[18666]  = 1;
  ram[18667]  = 1;
  ram[18668]  = 1;
  ram[18669]  = 1;
  ram[18670]  = 1;
  ram[18671]  = 1;
  ram[18672]  = 1;
  ram[18673]  = 1;
  ram[18674]  = 1;
  ram[18675]  = 1;
  ram[18676]  = 1;
  ram[18677]  = 1;
  ram[18678]  = 1;
  ram[18679]  = 1;
  ram[18680]  = 1;
  ram[18681]  = 1;
  ram[18682]  = 1;
  ram[18683]  = 1;
  ram[18684]  = 1;
  ram[18685]  = 1;
  ram[18686]  = 1;
  ram[18687]  = 1;
  ram[18688]  = 1;
  ram[18689]  = 1;
  ram[18690]  = 1;
  ram[18691]  = 1;
  ram[18692]  = 1;
  ram[18693]  = 1;
  ram[18694]  = 1;
  ram[18695]  = 1;
  ram[18696]  = 1;
  ram[18697]  = 0;
  ram[18698]  = 1;
  ram[18699]  = 1;
  ram[18700]  = 1;
  ram[18701]  = 1;
  ram[18702]  = 1;
  ram[18703]  = 1;
  ram[18704]  = 1;
  ram[18705]  = 1;
  ram[18706]  = 1;
  ram[18707]  = 1;
  ram[18708]  = 1;
  ram[18709]  = 1;
  ram[18710]  = 1;
  ram[18711]  = 1;
  ram[18712]  = 1;
  ram[18713]  = 1;
  ram[18714]  = 1;
  ram[18715]  = 1;
  ram[18716]  = 1;
  ram[18717]  = 1;
  ram[18718]  = 1;
  ram[18719]  = 1;
  ram[18720]  = 1;
  ram[18721]  = 1;
  ram[18722]  = 0;
  ram[18723]  = 0;
  ram[18724]  = 1;
  ram[18725]  = 0;
  ram[18726]  = 0;
  ram[18727]  = 0;
  ram[18728]  = 1;
  ram[18729]  = 1;
  ram[18730]  = 1;
  ram[18731]  = 1;
  ram[18732]  = 1;
  ram[18733]  = 1;
  ram[18734]  = 1;
  ram[18735]  = 1;
  ram[18736]  = 1;
  ram[18737]  = 1;
  ram[18738]  = 1;
  ram[18739]  = 1;
  ram[18740]  = 1;
  ram[18741]  = 1;
  ram[18742]  = 1;
  ram[18743]  = 1;
  ram[18744]  = 1;
  ram[18745]  = 1;
  ram[18746]  = 1;
  ram[18747]  = 1;
  ram[18748]  = 1;
  ram[18749]  = 1;
  ram[18750]  = 1;
  ram[18751]  = 1;
  ram[18752]  = 1;
  ram[18753]  = 1;
  ram[18754]  = 1;
  ram[18755]  = 1;
  ram[18756]  = 1;
  ram[18757]  = 1;
  ram[18758]  = 1;
  ram[18759]  = 1;
  ram[18760]  = 1;
  ram[18761]  = 1;
  ram[18762]  = 1;
  ram[18763]  = 1;
  ram[18764]  = 1;
  ram[18765]  = 1;
  ram[18766]  = 1;
  ram[18767]  = 1;
  ram[18768]  = 1;
  ram[18769]  = 1;
  ram[18770]  = 1;
  ram[18771]  = 1;
  ram[18772]  = 1;
  ram[18773]  = 1;
  ram[18774]  = 1;
  ram[18775]  = 1;
  ram[18776]  = 1;
  ram[18777]  = 1;
  ram[18778]  = 1;
  ram[18779]  = 1;
  ram[18780]  = 1;
  ram[18781]  = 1;
  ram[18782]  = 1;
  ram[18783]  = 1;
  ram[18784]  = 1;
  ram[18785]  = 1;
  ram[18786]  = 1;
  ram[18787]  = 1;
  ram[18788]  = 1;
  ram[18789]  = 1;
  ram[18790]  = 1;
  ram[18791]  = 1;
  ram[18792]  = 1;
  ram[18793]  = 1;
  ram[18794]  = 1;
  ram[18795]  = 1;
  ram[18796]  = 1;
  ram[18797]  = 1;
  ram[18798]  = 1;
  ram[18799]  = 1;
  ram[18800]  = 1;
  ram[18801]  = 1;
  ram[18802]  = 1;
  ram[18803]  = 1;
  ram[18804]  = 1;
  ram[18805]  = 1;
  ram[18806]  = 1;
  ram[18807]  = 1;
  ram[18808]  = 1;
  ram[18809]  = 1;
  ram[18810]  = 1;
  ram[18811]  = 1;
  ram[18812]  = 1;
  ram[18813]  = 1;
  ram[18814]  = 1;
  ram[18815]  = 1;
  ram[18816]  = 1;
  ram[18817]  = 1;
  ram[18818]  = 1;
  ram[18819]  = 1;
  ram[18820]  = 1;
  ram[18821]  = 1;
  ram[18822]  = 1;
  ram[18823]  = 1;
  ram[18824]  = 1;
  ram[18825]  = 1;
  ram[18826]  = 1;
  ram[18827]  = 1;
  ram[18828]  = 1;
  ram[18829]  = 1;
  ram[18830]  = 1;
  ram[18831]  = 1;
  ram[18832]  = 1;
  ram[18833]  = 1;
  ram[18834]  = 1;
  ram[18835]  = 1;
  ram[18836]  = 1;
  ram[18837]  = 1;
  ram[18838]  = 1;
  ram[18839]  = 1;
  ram[18840]  = 1;
  ram[18841]  = 1;
  ram[18842]  = 1;
  ram[18843]  = 1;
  ram[18844]  = 1;
  ram[18845]  = 1;
  ram[18846]  = 1;
  ram[18847]  = 1;
  ram[18848]  = 1;
  ram[18849]  = 1;
  ram[18850]  = 1;
  ram[18851]  = 1;
  ram[18852]  = 1;
  ram[18853]  = 1;
  ram[18854]  = 1;
  ram[18855]  = 1;
  ram[18856]  = 1;
  ram[18857]  = 1;
  ram[18858]  = 1;
  ram[18859]  = 1;
  ram[18860]  = 1;
  ram[18861]  = 1;
  ram[18862]  = 1;
  ram[18863]  = 1;
  ram[18864]  = 1;
  ram[18865]  = 1;
  ram[18866]  = 1;
  ram[18867]  = 1;
  ram[18868]  = 1;
  ram[18869]  = 1;
  ram[18870]  = 1;
  ram[18871]  = 1;
  ram[18872]  = 1;
  ram[18873]  = 1;
  ram[18874]  = 1;
  ram[18875]  = 1;
  ram[18876]  = 1;
  ram[18877]  = 1;
  ram[18878]  = 1;
  ram[18879]  = 1;
  ram[18880]  = 1;
  ram[18881]  = 1;
  ram[18882]  = 1;
  ram[18883]  = 1;
  ram[18884]  = 1;
  ram[18885]  = 1;
  ram[18886]  = 1;
  ram[18887]  = 1;
  ram[18888]  = 1;
  ram[18889]  = 1;
  ram[18890]  = 1;
  ram[18891]  = 1;
  ram[18892]  = 1;
  ram[18893]  = 1;
  ram[18894]  = 1;
  ram[18895]  = 1;
  ram[18896]  = 1;
  ram[18897]  = 1;
  ram[18898]  = 1;
  ram[18899]  = 1;
  ram[18900]  = 1;
  ram[18901]  = 1;
  ram[18902]  = 1;
  ram[18903]  = 1;
  ram[18904]  = 1;
  ram[18905]  = 1;
  ram[18906]  = 1;
  ram[18907]  = 1;
  ram[18908]  = 1;
  ram[18909]  = 1;
  ram[18910]  = 1;
  ram[18911]  = 1;
  ram[18912]  = 1;
  ram[18913]  = 1;
  ram[18914]  = 1;
  ram[18915]  = 1;
  ram[18916]  = 1;
  ram[18917]  = 1;
  ram[18918]  = 1;
  ram[18919]  = 1;
  ram[18920]  = 1;
  ram[18921]  = 1;
  ram[18922]  = 1;
  ram[18923]  = 1;
  ram[18924]  = 1;
  ram[18925]  = 1;
  ram[18926]  = 1;
  ram[18927]  = 1;
  ram[18928]  = 1;
  ram[18929]  = 1;
  ram[18930]  = 1;
  ram[18931]  = 1;
  ram[18932]  = 1;
  ram[18933]  = 1;
  ram[18934]  = 1;
  ram[18935]  = 1;
  ram[18936]  = 1;
  ram[18937]  = 1;
  ram[18938]  = 1;
  ram[18939]  = 1;
  ram[18940]  = 1;
  ram[18941]  = 1;
  ram[18942]  = 1;
  ram[18943]  = 1;
  ram[18944]  = 1;
  ram[18945]  = 0;
  ram[18946]  = 1;
  ram[18947]  = 1;
  ram[18948]  = 1;
  ram[18949]  = 1;
  ram[18950]  = 0;
  ram[18951]  = 0;
  ram[18952]  = 1;
  ram[18953]  = 1;
  ram[18954]  = 1;
  ram[18955]  = 1;
  ram[18956]  = 1;
  ram[18957]  = 1;
  ram[18958]  = 1;
  ram[18959]  = 1;
  ram[18960]  = 1;
  ram[18961]  = 1;
  ram[18962]  = 1;
  ram[18963]  = 1;
  ram[18964]  = 1;
  ram[18965]  = 1;
  ram[18966]  = 1;
  ram[18967]  = 1;
  ram[18968]  = 1;
  ram[18969]  = 1;
  ram[18970]  = 1;
  ram[18971]  = 1;
  ram[18972]  = 1;
  ram[18973]  = 1;
  ram[18974]  = 1;
  ram[18975]  = 1;
  ram[18976]  = 1;
  ram[18977]  = 1;
  ram[18978]  = 1;
  ram[18979]  = 1;
  ram[18980]  = 1;
  ram[18981]  = 1;
  ram[18982]  = 1;
  ram[18983]  = 1;
  ram[18984]  = 1;
  ram[18985]  = 1;
  ram[18986]  = 1;
  ram[18987]  = 1;
  ram[18988]  = 1;
  ram[18989]  = 1;
  ram[18990]  = 1;
  ram[18991]  = 0;
  ram[18992]  = 1;
  ram[18993]  = 1;
  ram[18994]  = 1;
  ram[18995]  = 1;
  ram[18996]  = 1;
  ram[18997]  = 0;
  ram[18998]  = 1;
  ram[18999]  = 1;
  ram[19000]  = 1;
  ram[19001]  = 1;
  ram[19002]  = 1;
  ram[19003]  = 1;
  ram[19004]  = 1;
  ram[19005]  = 1;
  ram[19006]  = 1;
  ram[19007]  = 1;
  ram[19008]  = 1;
  ram[19009]  = 1;
  ram[19010]  = 1;
  ram[19011]  = 1;
  ram[19012]  = 1;
  ram[19013]  = 1;
  ram[19014]  = 1;
  ram[19015]  = 1;
  ram[19016]  = 1;
  ram[19017]  = 1;
  ram[19018]  = 1;
  ram[19019]  = 1;
  ram[19020]  = 1;
  ram[19021]  = 1;
  ram[19022]  = 0;
  ram[19023]  = 1;
  ram[19024]  = 1;
  ram[19025]  = 1;
  ram[19026]  = 1;
  ram[19027]  = 0;
  ram[19028]  = 0;
  ram[19029]  = 1;
  ram[19030]  = 1;
  ram[19031]  = 1;
  ram[19032]  = 1;
  ram[19033]  = 1;
  ram[19034]  = 1;
  ram[19035]  = 1;
  ram[19036]  = 1;
  ram[19037]  = 1;
  ram[19038]  = 1;
  ram[19039]  = 1;
  ram[19040]  = 1;
  ram[19041]  = 1;
  ram[19042]  = 1;
  ram[19043]  = 1;
  ram[19044]  = 1;
  ram[19045]  = 1;
  ram[19046]  = 1;
  ram[19047]  = 1;
  ram[19048]  = 1;
  ram[19049]  = 1;
  ram[19050]  = 1;
  ram[19051]  = 1;
  ram[19052]  = 1;
  ram[19053]  = 1;
  ram[19054]  = 1;
  ram[19055]  = 1;
  ram[19056]  = 1;
  ram[19057]  = 1;
  ram[19058]  = 1;
  ram[19059]  = 1;
  ram[19060]  = 1;
  ram[19061]  = 1;
  ram[19062]  = 1;
  ram[19063]  = 1;
  ram[19064]  = 1;
  ram[19065]  = 1;
  ram[19066]  = 1;
  ram[19067]  = 1;
  ram[19068]  = 1;
  ram[19069]  = 1;
  ram[19070]  = 1;
  ram[19071]  = 1;
  ram[19072]  = 1;
  ram[19073]  = 1;
  ram[19074]  = 1;
  ram[19075]  = 1;
  ram[19076]  = 1;
  ram[19077]  = 1;
  ram[19078]  = 1;
  ram[19079]  = 1;
  ram[19080]  = 0;
  ram[19081]  = 1;
  ram[19082]  = 1;
  ram[19083]  = 1;
  ram[19084]  = 1;
  ram[19085]  = 1;
  ram[19086]  = 1;
  ram[19087]  = 1;
  ram[19088]  = 1;
  ram[19089]  = 1;
  ram[19090]  = 1;
  ram[19091]  = 1;
  ram[19092]  = 1;
  ram[19093]  = 1;
  ram[19094]  = 1;
  ram[19095]  = 1;
  ram[19096]  = 1;
  ram[19097]  = 1;
  ram[19098]  = 1;
  ram[19099]  = 1;
  ram[19100]  = 1;
  ram[19101]  = 1;
  ram[19102]  = 1;
  ram[19103]  = 1;
  ram[19104]  = 1;
  ram[19105]  = 1;
  ram[19106]  = 1;
  ram[19107]  = 1;
  ram[19108]  = 1;
  ram[19109]  = 1;
  ram[19110]  = 1;
  ram[19111]  = 1;
  ram[19112]  = 1;
  ram[19113]  = 1;
  ram[19114]  = 1;
  ram[19115]  = 1;
  ram[19116]  = 1;
  ram[19117]  = 1;
  ram[19118]  = 1;
  ram[19119]  = 1;
  ram[19120]  = 1;
  ram[19121]  = 1;
  ram[19122]  = 1;
  ram[19123]  = 1;
  ram[19124]  = 1;
  ram[19125]  = 0;
  ram[19126]  = 1;
  ram[19127]  = 1;
  ram[19128]  = 1;
  ram[19129]  = 1;
  ram[19130]  = 1;
  ram[19131]  = 1;
  ram[19132]  = 1;
  ram[19133]  = 1;
  ram[19134]  = 1;
  ram[19135]  = 1;
  ram[19136]  = 1;
  ram[19137]  = 1;
  ram[19138]  = 1;
  ram[19139]  = 1;
  ram[19140]  = 1;
  ram[19141]  = 1;
  ram[19142]  = 1;
  ram[19143]  = 1;
  ram[19144]  = 1;
  ram[19145]  = 1;
  ram[19146]  = 1;
  ram[19147]  = 0;
  ram[19148]  = 1;
  ram[19149]  = 1;
  ram[19150]  = 1;
  ram[19151]  = 1;
  ram[19152]  = 1;
  ram[19153]  = 1;
  ram[19154]  = 1;
  ram[19155]  = 1;
  ram[19156]  = 1;
  ram[19157]  = 1;
  ram[19158]  = 1;
  ram[19159]  = 1;
  ram[19160]  = 1;
  ram[19161]  = 1;
  ram[19162]  = 1;
  ram[19163]  = 1;
  ram[19164]  = 1;
  ram[19165]  = 1;
  ram[19166]  = 1;
  ram[19167]  = 1;
  ram[19168]  = 1;
  ram[19169]  = 1;
  ram[19170]  = 1;
  ram[19171]  = 1;
  ram[19172]  = 1;
  ram[19173]  = 1;
  ram[19174]  = 1;
  ram[19175]  = 1;
  ram[19176]  = 1;
  ram[19177]  = 1;
  ram[19178]  = 1;
  ram[19179]  = 1;
  ram[19180]  = 1;
  ram[19181]  = 1;
  ram[19182]  = 1;
  ram[19183]  = 1;
  ram[19184]  = 1;
  ram[19185]  = 1;
  ram[19186]  = 1;
  ram[19187]  = 1;
  ram[19188]  = 1;
  ram[19189]  = 1;
  ram[19190]  = 1;
  ram[19191]  = 1;
  ram[19192]  = 1;
  ram[19193]  = 1;
  ram[19194]  = 1;
  ram[19195]  = 1;
  ram[19196]  = 1;
  ram[19197]  = 1;
  ram[19198]  = 1;
  ram[19199]  = 1;
  ram[19200]  = 1;
  ram[19201]  = 1;
  ram[19202]  = 1;
  ram[19203]  = 1;
  ram[19204]  = 1;
  ram[19205]  = 1;
  ram[19206]  = 1;
  ram[19207]  = 1;
  ram[19208]  = 1;
  ram[19209]  = 1;
  ram[19210]  = 1;
  ram[19211]  = 1;
  ram[19212]  = 1;
  ram[19213]  = 1;
  ram[19214]  = 1;
  ram[19215]  = 1;
  ram[19216]  = 1;
  ram[19217]  = 1;
  ram[19218]  = 1;
  ram[19219]  = 1;
  ram[19220]  = 1;
  ram[19221]  = 1;
  ram[19222]  = 1;
  ram[19223]  = 1;
  ram[19224]  = 1;
  ram[19225]  = 1;
  ram[19226]  = 1;
  ram[19227]  = 1;
  ram[19228]  = 1;
  ram[19229]  = 1;
  ram[19230]  = 1;
  ram[19231]  = 1;
  ram[19232]  = 1;
  ram[19233]  = 1;
  ram[19234]  = 1;
  ram[19235]  = 1;
  ram[19236]  = 1;
  ram[19237]  = 1;
  ram[19238]  = 1;
  ram[19239]  = 1;
  ram[19240]  = 1;
  ram[19241]  = 1;
  ram[19242]  = 1;
  ram[19243]  = 1;
  ram[19244]  = 1;
  ram[19245]  = 0;
  ram[19246]  = 1;
  ram[19247]  = 1;
  ram[19248]  = 1;
  ram[19249]  = 1;
  ram[19250]  = 1;
  ram[19251]  = 0;
  ram[19252]  = 1;
  ram[19253]  = 1;
  ram[19254]  = 1;
  ram[19255]  = 1;
  ram[19256]  = 1;
  ram[19257]  = 1;
  ram[19258]  = 1;
  ram[19259]  = 1;
  ram[19260]  = 1;
  ram[19261]  = 1;
  ram[19262]  = 1;
  ram[19263]  = 1;
  ram[19264]  = 1;
  ram[19265]  = 1;
  ram[19266]  = 1;
  ram[19267]  = 1;
  ram[19268]  = 1;
  ram[19269]  = 1;
  ram[19270]  = 1;
  ram[19271]  = 1;
  ram[19272]  = 1;
  ram[19273]  = 1;
  ram[19274]  = 1;
  ram[19275]  = 1;
  ram[19276]  = 1;
  ram[19277]  = 1;
  ram[19278]  = 1;
  ram[19279]  = 1;
  ram[19280]  = 1;
  ram[19281]  = 1;
  ram[19282]  = 1;
  ram[19283]  = 1;
  ram[19284]  = 1;
  ram[19285]  = 1;
  ram[19286]  = 1;
  ram[19287]  = 1;
  ram[19288]  = 1;
  ram[19289]  = 1;
  ram[19290]  = 1;
  ram[19291]  = 0;
  ram[19292]  = 1;
  ram[19293]  = 1;
  ram[19294]  = 1;
  ram[19295]  = 1;
  ram[19296]  = 1;
  ram[19297]  = 0;
  ram[19298]  = 1;
  ram[19299]  = 1;
  ram[19300]  = 1;
  ram[19301]  = 1;
  ram[19302]  = 1;
  ram[19303]  = 1;
  ram[19304]  = 1;
  ram[19305]  = 1;
  ram[19306]  = 1;
  ram[19307]  = 1;
  ram[19308]  = 1;
  ram[19309]  = 1;
  ram[19310]  = 1;
  ram[19311]  = 1;
  ram[19312]  = 1;
  ram[19313]  = 1;
  ram[19314]  = 1;
  ram[19315]  = 1;
  ram[19316]  = 1;
  ram[19317]  = 1;
  ram[19318]  = 1;
  ram[19319]  = 1;
  ram[19320]  = 1;
  ram[19321]  = 1;
  ram[19322]  = 0;
  ram[19323]  = 1;
  ram[19324]  = 1;
  ram[19325]  = 1;
  ram[19326]  = 1;
  ram[19327]  = 1;
  ram[19328]  = 0;
  ram[19329]  = 1;
  ram[19330]  = 1;
  ram[19331]  = 1;
  ram[19332]  = 1;
  ram[19333]  = 1;
  ram[19334]  = 1;
  ram[19335]  = 1;
  ram[19336]  = 1;
  ram[19337]  = 1;
  ram[19338]  = 1;
  ram[19339]  = 1;
  ram[19340]  = 1;
  ram[19341]  = 1;
  ram[19342]  = 1;
  ram[19343]  = 0;
  ram[19344]  = 1;
  ram[19345]  = 1;
  ram[19346]  = 1;
  ram[19347]  = 1;
  ram[19348]  = 0;
  ram[19349]  = 1;
  ram[19350]  = 1;
  ram[19351]  = 1;
  ram[19352]  = 1;
  ram[19353]  = 1;
  ram[19354]  = 1;
  ram[19355]  = 1;
  ram[19356]  = 1;
  ram[19357]  = 1;
  ram[19358]  = 1;
  ram[19359]  = 1;
  ram[19360]  = 1;
  ram[19361]  = 1;
  ram[19362]  = 1;
  ram[19363]  = 1;
  ram[19364]  = 1;
  ram[19365]  = 1;
  ram[19366]  = 1;
  ram[19367]  = 1;
  ram[19368]  = 1;
  ram[19369]  = 1;
  ram[19370]  = 1;
  ram[19371]  = 1;
  ram[19372]  = 1;
  ram[19373]  = 1;
  ram[19374]  = 1;
  ram[19375]  = 1;
  ram[19376]  = 1;
  ram[19377]  = 1;
  ram[19378]  = 1;
  ram[19379]  = 1;
  ram[19380]  = 0;
  ram[19381]  = 1;
  ram[19382]  = 1;
  ram[19383]  = 1;
  ram[19384]  = 1;
  ram[19385]  = 1;
  ram[19386]  = 1;
  ram[19387]  = 1;
  ram[19388]  = 1;
  ram[19389]  = 1;
  ram[19390]  = 1;
  ram[19391]  = 1;
  ram[19392]  = 1;
  ram[19393]  = 1;
  ram[19394]  = 1;
  ram[19395]  = 1;
  ram[19396]  = 1;
  ram[19397]  = 1;
  ram[19398]  = 1;
  ram[19399]  = 1;
  ram[19400]  = 1;
  ram[19401]  = 1;
  ram[19402]  = 1;
  ram[19403]  = 1;
  ram[19404]  = 1;
  ram[19405]  = 1;
  ram[19406]  = 1;
  ram[19407]  = 1;
  ram[19408]  = 1;
  ram[19409]  = 1;
  ram[19410]  = 1;
  ram[19411]  = 1;
  ram[19412]  = 1;
  ram[19413]  = 1;
  ram[19414]  = 1;
  ram[19415]  = 1;
  ram[19416]  = 1;
  ram[19417]  = 1;
  ram[19418]  = 1;
  ram[19419]  = 1;
  ram[19420]  = 1;
  ram[19421]  = 1;
  ram[19422]  = 1;
  ram[19423]  = 1;
  ram[19424]  = 1;
  ram[19425]  = 0;
  ram[19426]  = 1;
  ram[19427]  = 1;
  ram[19428]  = 1;
  ram[19429]  = 1;
  ram[19430]  = 1;
  ram[19431]  = 1;
  ram[19432]  = 1;
  ram[19433]  = 1;
  ram[19434]  = 1;
  ram[19435]  = 1;
  ram[19436]  = 1;
  ram[19437]  = 1;
  ram[19438]  = 1;
  ram[19439]  = 1;
  ram[19440]  = 1;
  ram[19441]  = 1;
  ram[19442]  = 1;
  ram[19443]  = 1;
  ram[19444]  = 1;
  ram[19445]  = 1;
  ram[19446]  = 1;
  ram[19447]  = 0;
  ram[19448]  = 1;
  ram[19449]  = 1;
  ram[19450]  = 1;
  ram[19451]  = 1;
  ram[19452]  = 1;
  ram[19453]  = 1;
  ram[19454]  = 1;
  ram[19455]  = 1;
  ram[19456]  = 1;
  ram[19457]  = 1;
  ram[19458]  = 1;
  ram[19459]  = 1;
  ram[19460]  = 1;
  ram[19461]  = 1;
  ram[19462]  = 1;
  ram[19463]  = 1;
  ram[19464]  = 1;
  ram[19465]  = 1;
  ram[19466]  = 1;
  ram[19467]  = 1;
  ram[19468]  = 1;
  ram[19469]  = 1;
  ram[19470]  = 1;
  ram[19471]  = 1;
  ram[19472]  = 1;
  ram[19473]  = 1;
  ram[19474]  = 1;
  ram[19475]  = 1;
  ram[19476]  = 1;
  ram[19477]  = 1;
  ram[19478]  = 1;
  ram[19479]  = 1;
  ram[19480]  = 1;
  ram[19481]  = 1;
  ram[19482]  = 1;
  ram[19483]  = 1;
  ram[19484]  = 1;
  ram[19485]  = 1;
  ram[19486]  = 1;
  ram[19487]  = 1;
  ram[19488]  = 1;
  ram[19489]  = 1;
  ram[19490]  = 1;
  ram[19491]  = 1;
  ram[19492]  = 1;
  ram[19493]  = 1;
  ram[19494]  = 1;
  ram[19495]  = 1;
  ram[19496]  = 1;
  ram[19497]  = 1;
  ram[19498]  = 1;
  ram[19499]  = 1;
  ram[19500]  = 1;
  ram[19501]  = 1;
  ram[19502]  = 1;
  ram[19503]  = 1;
  ram[19504]  = 1;
  ram[19505]  = 1;
  ram[19506]  = 1;
  ram[19507]  = 1;
  ram[19508]  = 1;
  ram[19509]  = 1;
  ram[19510]  = 1;
  ram[19511]  = 1;
  ram[19512]  = 1;
  ram[19513]  = 1;
  ram[19514]  = 1;
  ram[19515]  = 1;
  ram[19516]  = 1;
  ram[19517]  = 1;
  ram[19518]  = 1;
  ram[19519]  = 1;
  ram[19520]  = 1;
  ram[19521]  = 1;
  ram[19522]  = 1;
  ram[19523]  = 1;
  ram[19524]  = 1;
  ram[19525]  = 1;
  ram[19526]  = 1;
  ram[19527]  = 1;
  ram[19528]  = 1;
  ram[19529]  = 1;
  ram[19530]  = 1;
  ram[19531]  = 1;
  ram[19532]  = 1;
  ram[19533]  = 1;
  ram[19534]  = 1;
  ram[19535]  = 1;
  ram[19536]  = 1;
  ram[19537]  = 1;
  ram[19538]  = 1;
  ram[19539]  = 1;
  ram[19540]  = 1;
  ram[19541]  = 1;
  ram[19542]  = 1;
  ram[19543]  = 1;
  ram[19544]  = 1;
  ram[19545]  = 0;
  ram[19546]  = 1;
  ram[19547]  = 1;
  ram[19548]  = 1;
  ram[19549]  = 1;
  ram[19550]  = 1;
  ram[19551]  = 0;
  ram[19552]  = 0;
  ram[19553]  = 1;
  ram[19554]  = 1;
  ram[19555]  = 1;
  ram[19556]  = 1;
  ram[19557]  = 1;
  ram[19558]  = 1;
  ram[19559]  = 1;
  ram[19560]  = 1;
  ram[19561]  = 1;
  ram[19562]  = 1;
  ram[19563]  = 1;
  ram[19564]  = 1;
  ram[19565]  = 1;
  ram[19566]  = 1;
  ram[19567]  = 1;
  ram[19568]  = 1;
  ram[19569]  = 1;
  ram[19570]  = 1;
  ram[19571]  = 1;
  ram[19572]  = 1;
  ram[19573]  = 1;
  ram[19574]  = 1;
  ram[19575]  = 1;
  ram[19576]  = 1;
  ram[19577]  = 1;
  ram[19578]  = 1;
  ram[19579]  = 1;
  ram[19580]  = 1;
  ram[19581]  = 1;
  ram[19582]  = 1;
  ram[19583]  = 1;
  ram[19584]  = 1;
  ram[19585]  = 1;
  ram[19586]  = 1;
  ram[19587]  = 1;
  ram[19588]  = 1;
  ram[19589]  = 1;
  ram[19590]  = 1;
  ram[19591]  = 0;
  ram[19592]  = 1;
  ram[19593]  = 1;
  ram[19594]  = 1;
  ram[19595]  = 1;
  ram[19596]  = 1;
  ram[19597]  = 0;
  ram[19598]  = 1;
  ram[19599]  = 1;
  ram[19600]  = 1;
  ram[19601]  = 1;
  ram[19602]  = 1;
  ram[19603]  = 1;
  ram[19604]  = 1;
  ram[19605]  = 1;
  ram[19606]  = 1;
  ram[19607]  = 1;
  ram[19608]  = 1;
  ram[19609]  = 1;
  ram[19610]  = 1;
  ram[19611]  = 1;
  ram[19612]  = 1;
  ram[19613]  = 1;
  ram[19614]  = 1;
  ram[19615]  = 1;
  ram[19616]  = 1;
  ram[19617]  = 1;
  ram[19618]  = 1;
  ram[19619]  = 1;
  ram[19620]  = 1;
  ram[19621]  = 1;
  ram[19622]  = 0;
  ram[19623]  = 1;
  ram[19624]  = 1;
  ram[19625]  = 1;
  ram[19626]  = 1;
  ram[19627]  = 1;
  ram[19628]  = 0;
  ram[19629]  = 1;
  ram[19630]  = 1;
  ram[19631]  = 1;
  ram[19632]  = 1;
  ram[19633]  = 1;
  ram[19634]  = 1;
  ram[19635]  = 1;
  ram[19636]  = 1;
  ram[19637]  = 1;
  ram[19638]  = 1;
  ram[19639]  = 1;
  ram[19640]  = 1;
  ram[19641]  = 1;
  ram[19642]  = 0;
  ram[19643]  = 0;
  ram[19644]  = 1;
  ram[19645]  = 1;
  ram[19646]  = 1;
  ram[19647]  = 1;
  ram[19648]  = 0;
  ram[19649]  = 1;
  ram[19650]  = 1;
  ram[19651]  = 1;
  ram[19652]  = 1;
  ram[19653]  = 1;
  ram[19654]  = 1;
  ram[19655]  = 1;
  ram[19656]  = 1;
  ram[19657]  = 1;
  ram[19658]  = 1;
  ram[19659]  = 1;
  ram[19660]  = 1;
  ram[19661]  = 1;
  ram[19662]  = 1;
  ram[19663]  = 1;
  ram[19664]  = 1;
  ram[19665]  = 1;
  ram[19666]  = 1;
  ram[19667]  = 1;
  ram[19668]  = 1;
  ram[19669]  = 1;
  ram[19670]  = 1;
  ram[19671]  = 1;
  ram[19672]  = 1;
  ram[19673]  = 1;
  ram[19674]  = 1;
  ram[19675]  = 1;
  ram[19676]  = 1;
  ram[19677]  = 1;
  ram[19678]  = 1;
  ram[19679]  = 1;
  ram[19680]  = 0;
  ram[19681]  = 1;
  ram[19682]  = 1;
  ram[19683]  = 1;
  ram[19684]  = 1;
  ram[19685]  = 1;
  ram[19686]  = 1;
  ram[19687]  = 1;
  ram[19688]  = 1;
  ram[19689]  = 1;
  ram[19690]  = 1;
  ram[19691]  = 1;
  ram[19692]  = 1;
  ram[19693]  = 1;
  ram[19694]  = 1;
  ram[19695]  = 1;
  ram[19696]  = 1;
  ram[19697]  = 1;
  ram[19698]  = 1;
  ram[19699]  = 1;
  ram[19700]  = 1;
  ram[19701]  = 1;
  ram[19702]  = 1;
  ram[19703]  = 1;
  ram[19704]  = 1;
  ram[19705]  = 1;
  ram[19706]  = 1;
  ram[19707]  = 1;
  ram[19708]  = 1;
  ram[19709]  = 1;
  ram[19710]  = 1;
  ram[19711]  = 1;
  ram[19712]  = 1;
  ram[19713]  = 1;
  ram[19714]  = 1;
  ram[19715]  = 1;
  ram[19716]  = 1;
  ram[19717]  = 1;
  ram[19718]  = 1;
  ram[19719]  = 1;
  ram[19720]  = 1;
  ram[19721]  = 1;
  ram[19722]  = 1;
  ram[19723]  = 1;
  ram[19724]  = 1;
  ram[19725]  = 0;
  ram[19726]  = 1;
  ram[19727]  = 1;
  ram[19728]  = 1;
  ram[19729]  = 1;
  ram[19730]  = 1;
  ram[19731]  = 1;
  ram[19732]  = 1;
  ram[19733]  = 1;
  ram[19734]  = 1;
  ram[19735]  = 1;
  ram[19736]  = 1;
  ram[19737]  = 1;
  ram[19738]  = 1;
  ram[19739]  = 1;
  ram[19740]  = 1;
  ram[19741]  = 1;
  ram[19742]  = 1;
  ram[19743]  = 1;
  ram[19744]  = 1;
  ram[19745]  = 1;
  ram[19746]  = 0;
  ram[19747]  = 0;
  ram[19748]  = 1;
  ram[19749]  = 1;
  ram[19750]  = 1;
  ram[19751]  = 1;
  ram[19752]  = 1;
  ram[19753]  = 1;
  ram[19754]  = 1;
  ram[19755]  = 1;
  ram[19756]  = 1;
  ram[19757]  = 1;
  ram[19758]  = 1;
  ram[19759]  = 1;
  ram[19760]  = 1;
  ram[19761]  = 1;
  ram[19762]  = 1;
  ram[19763]  = 1;
  ram[19764]  = 1;
  ram[19765]  = 1;
  ram[19766]  = 1;
  ram[19767]  = 1;
  ram[19768]  = 1;
  ram[19769]  = 1;
  ram[19770]  = 1;
  ram[19771]  = 1;
  ram[19772]  = 1;
  ram[19773]  = 1;
  ram[19774]  = 1;
  ram[19775]  = 1;
  ram[19776]  = 1;
  ram[19777]  = 1;
  ram[19778]  = 1;
  ram[19779]  = 1;
  ram[19780]  = 1;
  ram[19781]  = 1;
  ram[19782]  = 1;
  ram[19783]  = 1;
  ram[19784]  = 1;
  ram[19785]  = 1;
  ram[19786]  = 1;
  ram[19787]  = 1;
  ram[19788]  = 1;
  ram[19789]  = 1;
  ram[19790]  = 1;
  ram[19791]  = 1;
  ram[19792]  = 1;
  ram[19793]  = 1;
  ram[19794]  = 1;
  ram[19795]  = 1;
  ram[19796]  = 1;
  ram[19797]  = 1;
  ram[19798]  = 1;
  ram[19799]  = 1;
  ram[19800]  = 1;
  ram[19801]  = 1;
  ram[19802]  = 1;
  ram[19803]  = 1;
  ram[19804]  = 1;
  ram[19805]  = 1;
  ram[19806]  = 1;
  ram[19807]  = 1;
  ram[19808]  = 1;
  ram[19809]  = 1;
  ram[19810]  = 1;
  ram[19811]  = 1;
  ram[19812]  = 1;
  ram[19813]  = 1;
  ram[19814]  = 1;
  ram[19815]  = 1;
  ram[19816]  = 1;
  ram[19817]  = 1;
  ram[19818]  = 1;
  ram[19819]  = 1;
  ram[19820]  = 1;
  ram[19821]  = 1;
  ram[19822]  = 1;
  ram[19823]  = 1;
  ram[19824]  = 1;
  ram[19825]  = 1;
  ram[19826]  = 1;
  ram[19827]  = 1;
  ram[19828]  = 1;
  ram[19829]  = 1;
  ram[19830]  = 1;
  ram[19831]  = 1;
  ram[19832]  = 1;
  ram[19833]  = 1;
  ram[19834]  = 1;
  ram[19835]  = 1;
  ram[19836]  = 1;
  ram[19837]  = 1;
  ram[19838]  = 1;
  ram[19839]  = 1;
  ram[19840]  = 1;
  ram[19841]  = 1;
  ram[19842]  = 1;
  ram[19843]  = 1;
  ram[19844]  = 1;
  ram[19845]  = 0;
  ram[19846]  = 1;
  ram[19847]  = 1;
  ram[19848]  = 1;
  ram[19849]  = 1;
  ram[19850]  = 1;
  ram[19851]  = 0;
  ram[19852]  = 0;
  ram[19853]  = 1;
  ram[19854]  = 1;
  ram[19855]  = 1;
  ram[19856]  = 1;
  ram[19857]  = 1;
  ram[19858]  = 1;
  ram[19859]  = 1;
  ram[19860]  = 1;
  ram[19861]  = 1;
  ram[19862]  = 1;
  ram[19863]  = 1;
  ram[19864]  = 1;
  ram[19865]  = 1;
  ram[19866]  = 1;
  ram[19867]  = 1;
  ram[19868]  = 1;
  ram[19869]  = 1;
  ram[19870]  = 1;
  ram[19871]  = 1;
  ram[19872]  = 1;
  ram[19873]  = 1;
  ram[19874]  = 1;
  ram[19875]  = 1;
  ram[19876]  = 1;
  ram[19877]  = 1;
  ram[19878]  = 1;
  ram[19879]  = 1;
  ram[19880]  = 1;
  ram[19881]  = 1;
  ram[19882]  = 1;
  ram[19883]  = 1;
  ram[19884]  = 1;
  ram[19885]  = 1;
  ram[19886]  = 1;
  ram[19887]  = 1;
  ram[19888]  = 1;
  ram[19889]  = 1;
  ram[19890]  = 1;
  ram[19891]  = 0;
  ram[19892]  = 1;
  ram[19893]  = 1;
  ram[19894]  = 1;
  ram[19895]  = 1;
  ram[19896]  = 1;
  ram[19897]  = 0;
  ram[19898]  = 1;
  ram[19899]  = 1;
  ram[19900]  = 1;
  ram[19901]  = 1;
  ram[19902]  = 1;
  ram[19903]  = 1;
  ram[19904]  = 1;
  ram[19905]  = 1;
  ram[19906]  = 1;
  ram[19907]  = 1;
  ram[19908]  = 1;
  ram[19909]  = 1;
  ram[19910]  = 1;
  ram[19911]  = 1;
  ram[19912]  = 1;
  ram[19913]  = 1;
  ram[19914]  = 1;
  ram[19915]  = 1;
  ram[19916]  = 1;
  ram[19917]  = 1;
  ram[19918]  = 1;
  ram[19919]  = 1;
  ram[19920]  = 1;
  ram[19921]  = 1;
  ram[19922]  = 0;
  ram[19923]  = 1;
  ram[19924]  = 1;
  ram[19925]  = 1;
  ram[19926]  = 1;
  ram[19927]  = 1;
  ram[19928]  = 0;
  ram[19929]  = 1;
  ram[19930]  = 1;
  ram[19931]  = 1;
  ram[19932]  = 1;
  ram[19933]  = 1;
  ram[19934]  = 1;
  ram[19935]  = 1;
  ram[19936]  = 1;
  ram[19937]  = 1;
  ram[19938]  = 1;
  ram[19939]  = 1;
  ram[19940]  = 1;
  ram[19941]  = 1;
  ram[19942]  = 0;
  ram[19943]  = 0;
  ram[19944]  = 1;
  ram[19945]  = 1;
  ram[19946]  = 1;
  ram[19947]  = 1;
  ram[19948]  = 0;
  ram[19949]  = 1;
  ram[19950]  = 1;
  ram[19951]  = 1;
  ram[19952]  = 1;
  ram[19953]  = 1;
  ram[19954]  = 1;
  ram[19955]  = 1;
  ram[19956]  = 1;
  ram[19957]  = 1;
  ram[19958]  = 1;
  ram[19959]  = 1;
  ram[19960]  = 1;
  ram[19961]  = 1;
  ram[19962]  = 1;
  ram[19963]  = 1;
  ram[19964]  = 1;
  ram[19965]  = 1;
  ram[19966]  = 1;
  ram[19967]  = 1;
  ram[19968]  = 1;
  ram[19969]  = 1;
  ram[19970]  = 1;
  ram[19971]  = 1;
  ram[19972]  = 1;
  ram[19973]  = 1;
  ram[19974]  = 1;
  ram[19975]  = 1;
  ram[19976]  = 1;
  ram[19977]  = 1;
  ram[19978]  = 1;
  ram[19979]  = 1;
  ram[19980]  = 0;
  ram[19981]  = 1;
  ram[19982]  = 1;
  ram[19983]  = 1;
  ram[19984]  = 1;
  ram[19985]  = 1;
  ram[19986]  = 1;
  ram[19987]  = 1;
  ram[19988]  = 1;
  ram[19989]  = 1;
  ram[19990]  = 1;
  ram[19991]  = 1;
  ram[19992]  = 1;
  ram[19993]  = 1;
  ram[19994]  = 1;
  ram[19995]  = 1;
  ram[19996]  = 1;
  ram[19997]  = 1;
  ram[19998]  = 1;
  ram[19999]  = 1;
  ram[20000]  = 1;
  ram[20001]  = 1;
  ram[20002]  = 1;
  ram[20003]  = 1;
  ram[20004]  = 1;
  ram[20005]  = 1;
  ram[20006]  = 1;
  ram[20007]  = 1;
  ram[20008]  = 1;
  ram[20009]  = 1;
  ram[20010]  = 1;
  ram[20011]  = 1;
  ram[20012]  = 1;
  ram[20013]  = 1;
  ram[20014]  = 1;
  ram[20015]  = 1;
  ram[20016]  = 1;
  ram[20017]  = 1;
  ram[20018]  = 1;
  ram[20019]  = 1;
  ram[20020]  = 1;
  ram[20021]  = 1;
  ram[20022]  = 1;
  ram[20023]  = 1;
  ram[20024]  = 1;
  ram[20025]  = 0;
  ram[20026]  = 1;
  ram[20027]  = 1;
  ram[20028]  = 1;
  ram[20029]  = 1;
  ram[20030]  = 1;
  ram[20031]  = 1;
  ram[20032]  = 1;
  ram[20033]  = 1;
  ram[20034]  = 1;
  ram[20035]  = 1;
  ram[20036]  = 1;
  ram[20037]  = 1;
  ram[20038]  = 1;
  ram[20039]  = 1;
  ram[20040]  = 1;
  ram[20041]  = 1;
  ram[20042]  = 1;
  ram[20043]  = 1;
  ram[20044]  = 1;
  ram[20045]  = 1;
  ram[20046]  = 0;
  ram[20047]  = 0;
  ram[20048]  = 1;
  ram[20049]  = 1;
  ram[20050]  = 1;
  ram[20051]  = 1;
  ram[20052]  = 1;
  ram[20053]  = 1;
  ram[20054]  = 1;
  ram[20055]  = 1;
  ram[20056]  = 1;
  ram[20057]  = 1;
  ram[20058]  = 1;
  ram[20059]  = 1;
  ram[20060]  = 1;
  ram[20061]  = 1;
  ram[20062]  = 1;
  ram[20063]  = 1;
  ram[20064]  = 1;
  ram[20065]  = 1;
  ram[20066]  = 1;
  ram[20067]  = 1;
  ram[20068]  = 1;
  ram[20069]  = 1;
  ram[20070]  = 1;
  ram[20071]  = 1;
  ram[20072]  = 1;
  ram[20073]  = 1;
  ram[20074]  = 1;
  ram[20075]  = 1;
  ram[20076]  = 1;
  ram[20077]  = 1;
  ram[20078]  = 1;
  ram[20079]  = 1;
  ram[20080]  = 1;
  ram[20081]  = 1;
  ram[20082]  = 1;
  ram[20083]  = 1;
  ram[20084]  = 1;
  ram[20085]  = 1;
  ram[20086]  = 1;
  ram[20087]  = 1;
  ram[20088]  = 1;
  ram[20089]  = 1;
  ram[20090]  = 1;
  ram[20091]  = 1;
  ram[20092]  = 1;
  ram[20093]  = 1;
  ram[20094]  = 1;
  ram[20095]  = 1;
  ram[20096]  = 1;
  ram[20097]  = 1;
  ram[20098]  = 1;
  ram[20099]  = 1;
  ram[20100]  = 1;
  ram[20101]  = 1;
  ram[20102]  = 1;
  ram[20103]  = 1;
  ram[20104]  = 1;
  ram[20105]  = 1;
  ram[20106]  = 1;
  ram[20107]  = 1;
  ram[20108]  = 1;
  ram[20109]  = 1;
  ram[20110]  = 1;
  ram[20111]  = 1;
  ram[20112]  = 1;
  ram[20113]  = 1;
  ram[20114]  = 1;
  ram[20115]  = 1;
  ram[20116]  = 1;
  ram[20117]  = 1;
  ram[20118]  = 1;
  ram[20119]  = 1;
  ram[20120]  = 1;
  ram[20121]  = 1;
  ram[20122]  = 1;
  ram[20123]  = 1;
  ram[20124]  = 1;
  ram[20125]  = 1;
  ram[20126]  = 1;
  ram[20127]  = 1;
  ram[20128]  = 1;
  ram[20129]  = 1;
  ram[20130]  = 1;
  ram[20131]  = 1;
  ram[20132]  = 1;
  ram[20133]  = 1;
  ram[20134]  = 1;
  ram[20135]  = 1;
  ram[20136]  = 1;
  ram[20137]  = 1;
  ram[20138]  = 1;
  ram[20139]  = 1;
  ram[20140]  = 1;
  ram[20141]  = 1;
  ram[20142]  = 1;
  ram[20143]  = 1;
  ram[20144]  = 1;
  ram[20145]  = 0;
  ram[20146]  = 1;
  ram[20147]  = 1;
  ram[20148]  = 1;
  ram[20149]  = 1;
  ram[20150]  = 1;
  ram[20151]  = 0;
  ram[20152]  = 0;
  ram[20153]  = 1;
  ram[20154]  = 1;
  ram[20155]  = 0;
  ram[20156]  = 1;
  ram[20157]  = 0;
  ram[20158]  = 0;
  ram[20159]  = 0;
  ram[20160]  = 1;
  ram[20161]  = 1;
  ram[20162]  = 1;
  ram[20163]  = 0;
  ram[20164]  = 0;
  ram[20165]  = 0;
  ram[20166]  = 0;
  ram[20167]  = 1;
  ram[20168]  = 1;
  ram[20169]  = 1;
  ram[20170]  = 1;
  ram[20171]  = 0;
  ram[20172]  = 0;
  ram[20173]  = 0;
  ram[20174]  = 0;
  ram[20175]  = 1;
  ram[20176]  = 1;
  ram[20177]  = 1;
  ram[20178]  = 0;
  ram[20179]  = 0;
  ram[20180]  = 0;
  ram[20181]  = 0;
  ram[20182]  = 1;
  ram[20183]  = 1;
  ram[20184]  = 1;
  ram[20185]  = 1;
  ram[20186]  = 1;
  ram[20187]  = 1;
  ram[20188]  = 1;
  ram[20189]  = 1;
  ram[20190]  = 0;
  ram[20191]  = 0;
  ram[20192]  = 0;
  ram[20193]  = 0;
  ram[20194]  = 0;
  ram[20195]  = 1;
  ram[20196]  = 1;
  ram[20197]  = 0;
  ram[20198]  = 1;
  ram[20199]  = 0;
  ram[20200]  = 0;
  ram[20201]  = 0;
  ram[20202]  = 0;
  ram[20203]  = 1;
  ram[20204]  = 1;
  ram[20205]  = 1;
  ram[20206]  = 1;
  ram[20207]  = 1;
  ram[20208]  = 0;
  ram[20209]  = 0;
  ram[20210]  = 0;
  ram[20211]  = 0;
  ram[20212]  = 1;
  ram[20213]  = 1;
  ram[20214]  = 1;
  ram[20215]  = 1;
  ram[20216]  = 1;
  ram[20217]  = 1;
  ram[20218]  = 1;
  ram[20219]  = 1;
  ram[20220]  = 1;
  ram[20221]  = 1;
  ram[20222]  = 0;
  ram[20223]  = 1;
  ram[20224]  = 1;
  ram[20225]  = 1;
  ram[20226]  = 1;
  ram[20227]  = 1;
  ram[20228]  = 0;
  ram[20229]  = 1;
  ram[20230]  = 1;
  ram[20231]  = 1;
  ram[20232]  = 0;
  ram[20233]  = 1;
  ram[20234]  = 1;
  ram[20235]  = 1;
  ram[20236]  = 1;
  ram[20237]  = 1;
  ram[20238]  = 0;
  ram[20239]  = 1;
  ram[20240]  = 1;
  ram[20241]  = 0;
  ram[20242]  = 0;
  ram[20243]  = 0;
  ram[20244]  = 0;
  ram[20245]  = 0;
  ram[20246]  = 1;
  ram[20247]  = 0;
  ram[20248]  = 0;
  ram[20249]  = 0;
  ram[20250]  = 0;
  ram[20251]  = 0;
  ram[20252]  = 1;
  ram[20253]  = 1;
  ram[20254]  = 1;
  ram[20255]  = 0;
  ram[20256]  = 0;
  ram[20257]  = 0;
  ram[20258]  = 0;
  ram[20259]  = 0;
  ram[20260]  = 1;
  ram[20261]  = 1;
  ram[20262]  = 1;
  ram[20263]  = 1;
  ram[20264]  = 0;
  ram[20265]  = 0;
  ram[20266]  = 1;
  ram[20267]  = 0;
  ram[20268]  = 0;
  ram[20269]  = 0;
  ram[20270]  = 0;
  ram[20271]  = 1;
  ram[20272]  = 1;
  ram[20273]  = 1;
  ram[20274]  = 1;
  ram[20275]  = 1;
  ram[20276]  = 1;
  ram[20277]  = 1;
  ram[20278]  = 1;
  ram[20279]  = 0;
  ram[20280]  = 0;
  ram[20281]  = 0;
  ram[20282]  = 0;
  ram[20283]  = 0;
  ram[20284]  = 1;
  ram[20285]  = 1;
  ram[20286]  = 1;
  ram[20287]  = 0;
  ram[20288]  = 0;
  ram[20289]  = 0;
  ram[20290]  = 0;
  ram[20291]  = 0;
  ram[20292]  = 1;
  ram[20293]  = 1;
  ram[20294]  = 1;
  ram[20295]  = 1;
  ram[20296]  = 1;
  ram[20297]  = 1;
  ram[20298]  = 1;
  ram[20299]  = 1;
  ram[20300]  = 1;
  ram[20301]  = 0;
  ram[20302]  = 1;
  ram[20303]  = 1;
  ram[20304]  = 0;
  ram[20305]  = 0;
  ram[20306]  = 1;
  ram[20307]  = 1;
  ram[20308]  = 1;
  ram[20309]  = 0;
  ram[20310]  = 0;
  ram[20311]  = 0;
  ram[20312]  = 0;
  ram[20313]  = 1;
  ram[20314]  = 1;
  ram[20315]  = 1;
  ram[20316]  = 1;
  ram[20317]  = 0;
  ram[20318]  = 0;
  ram[20319]  = 0;
  ram[20320]  = 0;
  ram[20321]  = 0;
  ram[20322]  = 1;
  ram[20323]  = 1;
  ram[20324]  = 0;
  ram[20325]  = 0;
  ram[20326]  = 0;
  ram[20327]  = 0;
  ram[20328]  = 0;
  ram[20329]  = 1;
  ram[20330]  = 1;
  ram[20331]  = 0;
  ram[20332]  = 0;
  ram[20333]  = 0;
  ram[20334]  = 0;
  ram[20335]  = 0;
  ram[20336]  = 1;
  ram[20337]  = 1;
  ram[20338]  = 1;
  ram[20339]  = 1;
  ram[20340]  = 0;
  ram[20341]  = 1;
  ram[20342]  = 0;
  ram[20343]  = 0;
  ram[20344]  = 1;
  ram[20345]  = 0;
  ram[20346]  = 0;
  ram[20347]  = 0;
  ram[20348]  = 0;
  ram[20349]  = 0;
  ram[20350]  = 1;
  ram[20351]  = 1;
  ram[20352]  = 1;
  ram[20353]  = 1;
  ram[20354]  = 1;
  ram[20355]  = 1;
  ram[20356]  = 1;
  ram[20357]  = 1;
  ram[20358]  = 1;
  ram[20359]  = 1;
  ram[20360]  = 1;
  ram[20361]  = 1;
  ram[20362]  = 1;
  ram[20363]  = 1;
  ram[20364]  = 1;
  ram[20365]  = 1;
  ram[20366]  = 1;
  ram[20367]  = 1;
  ram[20368]  = 1;
  ram[20369]  = 1;
  ram[20370]  = 1;
  ram[20371]  = 1;
  ram[20372]  = 1;
  ram[20373]  = 1;
  ram[20374]  = 1;
  ram[20375]  = 1;
  ram[20376]  = 1;
  ram[20377]  = 1;
  ram[20378]  = 1;
  ram[20379]  = 1;
  ram[20380]  = 1;
  ram[20381]  = 1;
  ram[20382]  = 1;
  ram[20383]  = 1;
  ram[20384]  = 1;
  ram[20385]  = 1;
  ram[20386]  = 1;
  ram[20387]  = 1;
  ram[20388]  = 1;
  ram[20389]  = 1;
  ram[20390]  = 1;
  ram[20391]  = 1;
  ram[20392]  = 1;
  ram[20393]  = 1;
  ram[20394]  = 1;
  ram[20395]  = 1;
  ram[20396]  = 1;
  ram[20397]  = 1;
  ram[20398]  = 1;
  ram[20399]  = 1;
  ram[20400]  = 1;
  ram[20401]  = 1;
  ram[20402]  = 1;
  ram[20403]  = 1;
  ram[20404]  = 1;
  ram[20405]  = 1;
  ram[20406]  = 1;
  ram[20407]  = 1;
  ram[20408]  = 1;
  ram[20409]  = 1;
  ram[20410]  = 1;
  ram[20411]  = 1;
  ram[20412]  = 1;
  ram[20413]  = 1;
  ram[20414]  = 1;
  ram[20415]  = 1;
  ram[20416]  = 1;
  ram[20417]  = 1;
  ram[20418]  = 1;
  ram[20419]  = 1;
  ram[20420]  = 1;
  ram[20421]  = 1;
  ram[20422]  = 1;
  ram[20423]  = 1;
  ram[20424]  = 1;
  ram[20425]  = 1;
  ram[20426]  = 1;
  ram[20427]  = 1;
  ram[20428]  = 1;
  ram[20429]  = 1;
  ram[20430]  = 1;
  ram[20431]  = 1;
  ram[20432]  = 1;
  ram[20433]  = 1;
  ram[20434]  = 1;
  ram[20435]  = 1;
  ram[20436]  = 1;
  ram[20437]  = 1;
  ram[20438]  = 1;
  ram[20439]  = 1;
  ram[20440]  = 1;
  ram[20441]  = 1;
  ram[20442]  = 1;
  ram[20443]  = 1;
  ram[20444]  = 1;
  ram[20445]  = 0;
  ram[20446]  = 1;
  ram[20447]  = 1;
  ram[20448]  = 1;
  ram[20449]  = 1;
  ram[20450]  = 1;
  ram[20451]  = 0;
  ram[20452]  = 0;
  ram[20453]  = 1;
  ram[20454]  = 1;
  ram[20455]  = 0;
  ram[20456]  = 1;
  ram[20457]  = 0;
  ram[20458]  = 1;
  ram[20459]  = 1;
  ram[20460]  = 1;
  ram[20461]  = 1;
  ram[20462]  = 0;
  ram[20463]  = 0;
  ram[20464]  = 1;
  ram[20465]  = 1;
  ram[20466]  = 0;
  ram[20467]  = 1;
  ram[20468]  = 1;
  ram[20469]  = 1;
  ram[20470]  = 0;
  ram[20471]  = 0;
  ram[20472]  = 1;
  ram[20473]  = 1;
  ram[20474]  = 0;
  ram[20475]  = 0;
  ram[20476]  = 1;
  ram[20477]  = 1;
  ram[20478]  = 0;
  ram[20479]  = 1;
  ram[20480]  = 1;
  ram[20481]  = 1;
  ram[20482]  = 0;
  ram[20483]  = 1;
  ram[20484]  = 1;
  ram[20485]  = 1;
  ram[20486]  = 1;
  ram[20487]  = 1;
  ram[20488]  = 1;
  ram[20489]  = 1;
  ram[20490]  = 0;
  ram[20491]  = 0;
  ram[20492]  = 0;
  ram[20493]  = 0;
  ram[20494]  = 1;
  ram[20495]  = 1;
  ram[20496]  = 1;
  ram[20497]  = 0;
  ram[20498]  = 0;
  ram[20499]  = 0;
  ram[20500]  = 1;
  ram[20501]  = 0;
  ram[20502]  = 0;
  ram[20503]  = 1;
  ram[20504]  = 1;
  ram[20505]  = 1;
  ram[20506]  = 1;
  ram[20507]  = 1;
  ram[20508]  = 0;
  ram[20509]  = 1;
  ram[20510]  = 1;
  ram[20511]  = 0;
  ram[20512]  = 0;
  ram[20513]  = 1;
  ram[20514]  = 1;
  ram[20515]  = 1;
  ram[20516]  = 1;
  ram[20517]  = 1;
  ram[20518]  = 1;
  ram[20519]  = 1;
  ram[20520]  = 1;
  ram[20521]  = 1;
  ram[20522]  = 0;
  ram[20523]  = 1;
  ram[20524]  = 1;
  ram[20525]  = 1;
  ram[20526]  = 1;
  ram[20527]  = 0;
  ram[20528]  = 0;
  ram[20529]  = 1;
  ram[20530]  = 1;
  ram[20531]  = 1;
  ram[20532]  = 0;
  ram[20533]  = 1;
  ram[20534]  = 1;
  ram[20535]  = 1;
  ram[20536]  = 1;
  ram[20537]  = 1;
  ram[20538]  = 0;
  ram[20539]  = 1;
  ram[20540]  = 1;
  ram[20541]  = 0;
  ram[20542]  = 0;
  ram[20543]  = 0;
  ram[20544]  = 0;
  ram[20545]  = 0;
  ram[20546]  = 1;
  ram[20547]  = 0;
  ram[20548]  = 0;
  ram[20549]  = 0;
  ram[20550]  = 0;
  ram[20551]  = 0;
  ram[20552]  = 1;
  ram[20553]  = 1;
  ram[20554]  = 1;
  ram[20555]  = 0;
  ram[20556]  = 0;
  ram[20557]  = 1;
  ram[20558]  = 1;
  ram[20559]  = 0;
  ram[20560]  = 0;
  ram[20561]  = 1;
  ram[20562]  = 1;
  ram[20563]  = 1;
  ram[20564]  = 0;
  ram[20565]  = 0;
  ram[20566]  = 0;
  ram[20567]  = 0;
  ram[20568]  = 1;
  ram[20569]  = 0;
  ram[20570]  = 0;
  ram[20571]  = 1;
  ram[20572]  = 1;
  ram[20573]  = 1;
  ram[20574]  = 1;
  ram[20575]  = 1;
  ram[20576]  = 1;
  ram[20577]  = 1;
  ram[20578]  = 1;
  ram[20579]  = 0;
  ram[20580]  = 0;
  ram[20581]  = 0;
  ram[20582]  = 0;
  ram[20583]  = 1;
  ram[20584]  = 1;
  ram[20585]  = 1;
  ram[20586]  = 0;
  ram[20587]  = 0;
  ram[20588]  = 0;
  ram[20589]  = 1;
  ram[20590]  = 1;
  ram[20591]  = 0;
  ram[20592]  = 0;
  ram[20593]  = 1;
  ram[20594]  = 1;
  ram[20595]  = 1;
  ram[20596]  = 1;
  ram[20597]  = 1;
  ram[20598]  = 1;
  ram[20599]  = 1;
  ram[20600]  = 1;
  ram[20601]  = 0;
  ram[20602]  = 1;
  ram[20603]  = 0;
  ram[20604]  = 1;
  ram[20605]  = 1;
  ram[20606]  = 1;
  ram[20607]  = 1;
  ram[20608]  = 0;
  ram[20609]  = 0;
  ram[20610]  = 1;
  ram[20611]  = 1;
  ram[20612]  = 0;
  ram[20613]  = 0;
  ram[20614]  = 1;
  ram[20615]  = 1;
  ram[20616]  = 1;
  ram[20617]  = 0;
  ram[20618]  = 1;
  ram[20619]  = 1;
  ram[20620]  = 1;
  ram[20621]  = 0;
  ram[20622]  = 1;
  ram[20623]  = 1;
  ram[20624]  = 0;
  ram[20625]  = 0;
  ram[20626]  = 0;
  ram[20627]  = 0;
  ram[20628]  = 1;
  ram[20629]  = 1;
  ram[20630]  = 1;
  ram[20631]  = 0;
  ram[20632]  = 0;
  ram[20633]  = 1;
  ram[20634]  = 1;
  ram[20635]  = 0;
  ram[20636]  = 1;
  ram[20637]  = 1;
  ram[20638]  = 1;
  ram[20639]  = 1;
  ram[20640]  = 0;
  ram[20641]  = 1;
  ram[20642]  = 0;
  ram[20643]  = 1;
  ram[20644]  = 1;
  ram[20645]  = 0;
  ram[20646]  = 0;
  ram[20647]  = 0;
  ram[20648]  = 0;
  ram[20649]  = 0;
  ram[20650]  = 1;
  ram[20651]  = 1;
  ram[20652]  = 1;
  ram[20653]  = 1;
  ram[20654]  = 1;
  ram[20655]  = 1;
  ram[20656]  = 1;
  ram[20657]  = 1;
  ram[20658]  = 1;
  ram[20659]  = 1;
  ram[20660]  = 1;
  ram[20661]  = 1;
  ram[20662]  = 1;
  ram[20663]  = 1;
  ram[20664]  = 1;
  ram[20665]  = 1;
  ram[20666]  = 1;
  ram[20667]  = 1;
  ram[20668]  = 1;
  ram[20669]  = 1;
  ram[20670]  = 1;
  ram[20671]  = 1;
  ram[20672]  = 1;
  ram[20673]  = 1;
  ram[20674]  = 1;
  ram[20675]  = 1;
  ram[20676]  = 1;
  ram[20677]  = 1;
  ram[20678]  = 1;
  ram[20679]  = 1;
  ram[20680]  = 1;
  ram[20681]  = 1;
  ram[20682]  = 1;
  ram[20683]  = 1;
  ram[20684]  = 1;
  ram[20685]  = 1;
  ram[20686]  = 1;
  ram[20687]  = 1;
  ram[20688]  = 1;
  ram[20689]  = 1;
  ram[20690]  = 1;
  ram[20691]  = 1;
  ram[20692]  = 1;
  ram[20693]  = 1;
  ram[20694]  = 1;
  ram[20695]  = 1;
  ram[20696]  = 1;
  ram[20697]  = 1;
  ram[20698]  = 1;
  ram[20699]  = 1;
  ram[20700]  = 1;
  ram[20701]  = 1;
  ram[20702]  = 1;
  ram[20703]  = 1;
  ram[20704]  = 1;
  ram[20705]  = 1;
  ram[20706]  = 1;
  ram[20707]  = 1;
  ram[20708]  = 1;
  ram[20709]  = 1;
  ram[20710]  = 1;
  ram[20711]  = 1;
  ram[20712]  = 1;
  ram[20713]  = 1;
  ram[20714]  = 1;
  ram[20715]  = 1;
  ram[20716]  = 1;
  ram[20717]  = 1;
  ram[20718]  = 1;
  ram[20719]  = 1;
  ram[20720]  = 1;
  ram[20721]  = 1;
  ram[20722]  = 1;
  ram[20723]  = 1;
  ram[20724]  = 1;
  ram[20725]  = 1;
  ram[20726]  = 1;
  ram[20727]  = 1;
  ram[20728]  = 1;
  ram[20729]  = 1;
  ram[20730]  = 1;
  ram[20731]  = 1;
  ram[20732]  = 1;
  ram[20733]  = 1;
  ram[20734]  = 1;
  ram[20735]  = 1;
  ram[20736]  = 1;
  ram[20737]  = 1;
  ram[20738]  = 1;
  ram[20739]  = 1;
  ram[20740]  = 1;
  ram[20741]  = 1;
  ram[20742]  = 1;
  ram[20743]  = 1;
  ram[20744]  = 1;
  ram[20745]  = 0;
  ram[20746]  = 1;
  ram[20747]  = 1;
  ram[20748]  = 1;
  ram[20749]  = 1;
  ram[20750]  = 1;
  ram[20751]  = 0;
  ram[20752]  = 0;
  ram[20753]  = 1;
  ram[20754]  = 1;
  ram[20755]  = 0;
  ram[20756]  = 0;
  ram[20757]  = 1;
  ram[20758]  = 1;
  ram[20759]  = 1;
  ram[20760]  = 1;
  ram[20761]  = 0;
  ram[20762]  = 0;
  ram[20763]  = 1;
  ram[20764]  = 1;
  ram[20765]  = 1;
  ram[20766]  = 0;
  ram[20767]  = 0;
  ram[20768]  = 1;
  ram[20769]  = 1;
  ram[20770]  = 0;
  ram[20771]  = 1;
  ram[20772]  = 1;
  ram[20773]  = 1;
  ram[20774]  = 1;
  ram[20775]  = 0;
  ram[20776]  = 1;
  ram[20777]  = 1;
  ram[20778]  = 0;
  ram[20779]  = 1;
  ram[20780]  = 1;
  ram[20781]  = 1;
  ram[20782]  = 0;
  ram[20783]  = 1;
  ram[20784]  = 1;
  ram[20785]  = 1;
  ram[20786]  = 1;
  ram[20787]  = 1;
  ram[20788]  = 1;
  ram[20789]  = 1;
  ram[20790]  = 1;
  ram[20791]  = 0;
  ram[20792]  = 1;
  ram[20793]  = 1;
  ram[20794]  = 1;
  ram[20795]  = 1;
  ram[20796]  = 1;
  ram[20797]  = 0;
  ram[20798]  = 0;
  ram[20799]  = 1;
  ram[20800]  = 1;
  ram[20801]  = 1;
  ram[20802]  = 0;
  ram[20803]  = 0;
  ram[20804]  = 1;
  ram[20805]  = 1;
  ram[20806]  = 1;
  ram[20807]  = 0;
  ram[20808]  = 1;
  ram[20809]  = 1;
  ram[20810]  = 1;
  ram[20811]  = 1;
  ram[20812]  = 0;
  ram[20813]  = 0;
  ram[20814]  = 1;
  ram[20815]  = 1;
  ram[20816]  = 1;
  ram[20817]  = 1;
  ram[20818]  = 1;
  ram[20819]  = 1;
  ram[20820]  = 1;
  ram[20821]  = 1;
  ram[20822]  = 0;
  ram[20823]  = 1;
  ram[20824]  = 1;
  ram[20825]  = 1;
  ram[20826]  = 1;
  ram[20827]  = 0;
  ram[20828]  = 1;
  ram[20829]  = 1;
  ram[20830]  = 1;
  ram[20831]  = 1;
  ram[20832]  = 0;
  ram[20833]  = 1;
  ram[20834]  = 1;
  ram[20835]  = 1;
  ram[20836]  = 1;
  ram[20837]  = 1;
  ram[20838]  = 0;
  ram[20839]  = 1;
  ram[20840]  = 1;
  ram[20841]  = 1;
  ram[20842]  = 0;
  ram[20843]  = 0;
  ram[20844]  = 1;
  ram[20845]  = 1;
  ram[20846]  = 1;
  ram[20847]  = 1;
  ram[20848]  = 0;
  ram[20849]  = 1;
  ram[20850]  = 1;
  ram[20851]  = 1;
  ram[20852]  = 1;
  ram[20853]  = 1;
  ram[20854]  = 0;
  ram[20855]  = 0;
  ram[20856]  = 1;
  ram[20857]  = 1;
  ram[20858]  = 1;
  ram[20859]  = 1;
  ram[20860]  = 0;
  ram[20861]  = 1;
  ram[20862]  = 1;
  ram[20863]  = 1;
  ram[20864]  = 0;
  ram[20865]  = 0;
  ram[20866]  = 0;
  ram[20867]  = 1;
  ram[20868]  = 1;
  ram[20869]  = 1;
  ram[20870]  = 0;
  ram[20871]  = 0;
  ram[20872]  = 1;
  ram[20873]  = 1;
  ram[20874]  = 1;
  ram[20875]  = 1;
  ram[20876]  = 1;
  ram[20877]  = 1;
  ram[20878]  = 1;
  ram[20879]  = 1;
  ram[20880]  = 0;
  ram[20881]  = 1;
  ram[20882]  = 1;
  ram[20883]  = 1;
  ram[20884]  = 1;
  ram[20885]  = 1;
  ram[20886]  = 0;
  ram[20887]  = 1;
  ram[20888]  = 1;
  ram[20889]  = 1;
  ram[20890]  = 1;
  ram[20891]  = 1;
  ram[20892]  = 0;
  ram[20893]  = 1;
  ram[20894]  = 1;
  ram[20895]  = 1;
  ram[20896]  = 1;
  ram[20897]  = 1;
  ram[20898]  = 1;
  ram[20899]  = 1;
  ram[20900]  = 1;
  ram[20901]  = 0;
  ram[20902]  = 0;
  ram[20903]  = 1;
  ram[20904]  = 1;
  ram[20905]  = 1;
  ram[20906]  = 1;
  ram[20907]  = 1;
  ram[20908]  = 0;
  ram[20909]  = 1;
  ram[20910]  = 1;
  ram[20911]  = 1;
  ram[20912]  = 1;
  ram[20913]  = 0;
  ram[20914]  = 1;
  ram[20915]  = 1;
  ram[20916]  = 1;
  ram[20917]  = 0;
  ram[20918]  = 1;
  ram[20919]  = 1;
  ram[20920]  = 1;
  ram[20921]  = 0;
  ram[20922]  = 1;
  ram[20923]  = 1;
  ram[20924]  = 1;
  ram[20925]  = 0;
  ram[20926]  = 1;
  ram[20927]  = 1;
  ram[20928]  = 1;
  ram[20929]  = 1;
  ram[20930]  = 0;
  ram[20931]  = 0;
  ram[20932]  = 1;
  ram[20933]  = 1;
  ram[20934]  = 1;
  ram[20935]  = 0;
  ram[20936]  = 0;
  ram[20937]  = 1;
  ram[20938]  = 1;
  ram[20939]  = 1;
  ram[20940]  = 0;
  ram[20941]  = 0;
  ram[20942]  = 1;
  ram[20943]  = 1;
  ram[20944]  = 1;
  ram[20945]  = 1;
  ram[20946]  = 0;
  ram[20947]  = 0;
  ram[20948]  = 1;
  ram[20949]  = 1;
  ram[20950]  = 1;
  ram[20951]  = 1;
  ram[20952]  = 1;
  ram[20953]  = 1;
  ram[20954]  = 1;
  ram[20955]  = 1;
  ram[20956]  = 1;
  ram[20957]  = 1;
  ram[20958]  = 1;
  ram[20959]  = 1;
  ram[20960]  = 1;
  ram[20961]  = 1;
  ram[20962]  = 1;
  ram[20963]  = 1;
  ram[20964]  = 1;
  ram[20965]  = 1;
  ram[20966]  = 1;
  ram[20967]  = 1;
  ram[20968]  = 1;
  ram[20969]  = 1;
  ram[20970]  = 1;
  ram[20971]  = 1;
  ram[20972]  = 1;
  ram[20973]  = 1;
  ram[20974]  = 1;
  ram[20975]  = 1;
  ram[20976]  = 1;
  ram[20977]  = 1;
  ram[20978]  = 1;
  ram[20979]  = 1;
  ram[20980]  = 1;
  ram[20981]  = 1;
  ram[20982]  = 1;
  ram[20983]  = 1;
  ram[20984]  = 1;
  ram[20985]  = 1;
  ram[20986]  = 1;
  ram[20987]  = 1;
  ram[20988]  = 1;
  ram[20989]  = 1;
  ram[20990]  = 1;
  ram[20991]  = 1;
  ram[20992]  = 1;
  ram[20993]  = 1;
  ram[20994]  = 1;
  ram[20995]  = 1;
  ram[20996]  = 1;
  ram[20997]  = 1;
  ram[20998]  = 1;
  ram[20999]  = 1;
  ram[21000]  = 1;
  ram[21001]  = 1;
  ram[21002]  = 1;
  ram[21003]  = 1;
  ram[21004]  = 1;
  ram[21005]  = 1;
  ram[21006]  = 1;
  ram[21007]  = 1;
  ram[21008]  = 1;
  ram[21009]  = 1;
  ram[21010]  = 1;
  ram[21011]  = 1;
  ram[21012]  = 1;
  ram[21013]  = 1;
  ram[21014]  = 1;
  ram[21015]  = 1;
  ram[21016]  = 1;
  ram[21017]  = 1;
  ram[21018]  = 1;
  ram[21019]  = 1;
  ram[21020]  = 1;
  ram[21021]  = 1;
  ram[21022]  = 1;
  ram[21023]  = 1;
  ram[21024]  = 1;
  ram[21025]  = 1;
  ram[21026]  = 1;
  ram[21027]  = 1;
  ram[21028]  = 1;
  ram[21029]  = 1;
  ram[21030]  = 1;
  ram[21031]  = 1;
  ram[21032]  = 1;
  ram[21033]  = 1;
  ram[21034]  = 1;
  ram[21035]  = 1;
  ram[21036]  = 1;
  ram[21037]  = 1;
  ram[21038]  = 1;
  ram[21039]  = 1;
  ram[21040]  = 1;
  ram[21041]  = 1;
  ram[21042]  = 1;
  ram[21043]  = 1;
  ram[21044]  = 1;
  ram[21045]  = 0;
  ram[21046]  = 1;
  ram[21047]  = 1;
  ram[21048]  = 1;
  ram[21049]  = 1;
  ram[21050]  = 1;
  ram[21051]  = 0;
  ram[21052]  = 1;
  ram[21053]  = 1;
  ram[21054]  = 1;
  ram[21055]  = 0;
  ram[21056]  = 0;
  ram[21057]  = 1;
  ram[21058]  = 1;
  ram[21059]  = 1;
  ram[21060]  = 1;
  ram[21061]  = 0;
  ram[21062]  = 1;
  ram[21063]  = 1;
  ram[21064]  = 1;
  ram[21065]  = 1;
  ram[21066]  = 1;
  ram[21067]  = 0;
  ram[21068]  = 1;
  ram[21069]  = 1;
  ram[21070]  = 0;
  ram[21071]  = 1;
  ram[21072]  = 1;
  ram[21073]  = 1;
  ram[21074]  = 1;
  ram[21075]  = 1;
  ram[21076]  = 1;
  ram[21077]  = 0;
  ram[21078]  = 0;
  ram[21079]  = 1;
  ram[21080]  = 1;
  ram[21081]  = 1;
  ram[21082]  = 1;
  ram[21083]  = 1;
  ram[21084]  = 1;
  ram[21085]  = 1;
  ram[21086]  = 1;
  ram[21087]  = 1;
  ram[21088]  = 1;
  ram[21089]  = 1;
  ram[21090]  = 1;
  ram[21091]  = 0;
  ram[21092]  = 1;
  ram[21093]  = 1;
  ram[21094]  = 1;
  ram[21095]  = 1;
  ram[21096]  = 1;
  ram[21097]  = 0;
  ram[21098]  = 1;
  ram[21099]  = 1;
  ram[21100]  = 1;
  ram[21101]  = 1;
  ram[21102]  = 1;
  ram[21103]  = 0;
  ram[21104]  = 1;
  ram[21105]  = 1;
  ram[21106]  = 1;
  ram[21107]  = 0;
  ram[21108]  = 1;
  ram[21109]  = 1;
  ram[21110]  = 1;
  ram[21111]  = 1;
  ram[21112]  = 1;
  ram[21113]  = 0;
  ram[21114]  = 1;
  ram[21115]  = 1;
  ram[21116]  = 1;
  ram[21117]  = 1;
  ram[21118]  = 1;
  ram[21119]  = 1;
  ram[21120]  = 1;
  ram[21121]  = 1;
  ram[21122]  = 0;
  ram[21123]  = 1;
  ram[21124]  = 1;
  ram[21125]  = 1;
  ram[21126]  = 0;
  ram[21127]  = 0;
  ram[21128]  = 1;
  ram[21129]  = 1;
  ram[21130]  = 1;
  ram[21131]  = 1;
  ram[21132]  = 0;
  ram[21133]  = 1;
  ram[21134]  = 1;
  ram[21135]  = 1;
  ram[21136]  = 1;
  ram[21137]  = 1;
  ram[21138]  = 0;
  ram[21139]  = 1;
  ram[21140]  = 1;
  ram[21141]  = 1;
  ram[21142]  = 0;
  ram[21143]  = 0;
  ram[21144]  = 1;
  ram[21145]  = 1;
  ram[21146]  = 1;
  ram[21147]  = 1;
  ram[21148]  = 0;
  ram[21149]  = 1;
  ram[21150]  = 1;
  ram[21151]  = 1;
  ram[21152]  = 1;
  ram[21153]  = 1;
  ram[21154]  = 0;
  ram[21155]  = 1;
  ram[21156]  = 1;
  ram[21157]  = 1;
  ram[21158]  = 1;
  ram[21159]  = 1;
  ram[21160]  = 0;
  ram[21161]  = 0;
  ram[21162]  = 1;
  ram[21163]  = 1;
  ram[21164]  = 0;
  ram[21165]  = 0;
  ram[21166]  = 1;
  ram[21167]  = 1;
  ram[21168]  = 1;
  ram[21169]  = 1;
  ram[21170]  = 0;
  ram[21171]  = 0;
  ram[21172]  = 1;
  ram[21173]  = 1;
  ram[21174]  = 1;
  ram[21175]  = 1;
  ram[21176]  = 1;
  ram[21177]  = 1;
  ram[21178]  = 1;
  ram[21179]  = 1;
  ram[21180]  = 0;
  ram[21181]  = 1;
  ram[21182]  = 1;
  ram[21183]  = 1;
  ram[21184]  = 1;
  ram[21185]  = 1;
  ram[21186]  = 0;
  ram[21187]  = 1;
  ram[21188]  = 1;
  ram[21189]  = 1;
  ram[21190]  = 1;
  ram[21191]  = 1;
  ram[21192]  = 0;
  ram[21193]  = 1;
  ram[21194]  = 1;
  ram[21195]  = 1;
  ram[21196]  = 1;
  ram[21197]  = 1;
  ram[21198]  = 1;
  ram[21199]  = 1;
  ram[21200]  = 1;
  ram[21201]  = 0;
  ram[21202]  = 0;
  ram[21203]  = 1;
  ram[21204]  = 1;
  ram[21205]  = 1;
  ram[21206]  = 1;
  ram[21207]  = 0;
  ram[21208]  = 0;
  ram[21209]  = 1;
  ram[21210]  = 1;
  ram[21211]  = 1;
  ram[21212]  = 1;
  ram[21213]  = 0;
  ram[21214]  = 0;
  ram[21215]  = 1;
  ram[21216]  = 0;
  ram[21217]  = 0;
  ram[21218]  = 1;
  ram[21219]  = 1;
  ram[21220]  = 1;
  ram[21221]  = 1;
  ram[21222]  = 1;
  ram[21223]  = 1;
  ram[21224]  = 1;
  ram[21225]  = 0;
  ram[21226]  = 1;
  ram[21227]  = 1;
  ram[21228]  = 1;
  ram[21229]  = 1;
  ram[21230]  = 1;
  ram[21231]  = 1;
  ram[21232]  = 1;
  ram[21233]  = 1;
  ram[21234]  = 1;
  ram[21235]  = 1;
  ram[21236]  = 0;
  ram[21237]  = 1;
  ram[21238]  = 1;
  ram[21239]  = 1;
  ram[21240]  = 0;
  ram[21241]  = 0;
  ram[21242]  = 1;
  ram[21243]  = 1;
  ram[21244]  = 1;
  ram[21245]  = 1;
  ram[21246]  = 0;
  ram[21247]  = 0;
  ram[21248]  = 1;
  ram[21249]  = 1;
  ram[21250]  = 1;
  ram[21251]  = 1;
  ram[21252]  = 1;
  ram[21253]  = 1;
  ram[21254]  = 1;
  ram[21255]  = 1;
  ram[21256]  = 1;
  ram[21257]  = 1;
  ram[21258]  = 1;
  ram[21259]  = 1;
  ram[21260]  = 1;
  ram[21261]  = 1;
  ram[21262]  = 1;
  ram[21263]  = 1;
  ram[21264]  = 1;
  ram[21265]  = 1;
  ram[21266]  = 1;
  ram[21267]  = 1;
  ram[21268]  = 1;
  ram[21269]  = 1;
  ram[21270]  = 1;
  ram[21271]  = 1;
  ram[21272]  = 1;
  ram[21273]  = 1;
  ram[21274]  = 1;
  ram[21275]  = 1;
  ram[21276]  = 1;
  ram[21277]  = 1;
  ram[21278]  = 1;
  ram[21279]  = 1;
  ram[21280]  = 1;
  ram[21281]  = 1;
  ram[21282]  = 1;
  ram[21283]  = 1;
  ram[21284]  = 1;
  ram[21285]  = 1;
  ram[21286]  = 1;
  ram[21287]  = 1;
  ram[21288]  = 1;
  ram[21289]  = 1;
  ram[21290]  = 1;
  ram[21291]  = 1;
  ram[21292]  = 1;
  ram[21293]  = 1;
  ram[21294]  = 1;
  ram[21295]  = 1;
  ram[21296]  = 1;
  ram[21297]  = 1;
  ram[21298]  = 1;
  ram[21299]  = 1;
  ram[21300]  = 1;
  ram[21301]  = 1;
  ram[21302]  = 1;
  ram[21303]  = 1;
  ram[21304]  = 1;
  ram[21305]  = 1;
  ram[21306]  = 1;
  ram[21307]  = 1;
  ram[21308]  = 1;
  ram[21309]  = 1;
  ram[21310]  = 1;
  ram[21311]  = 1;
  ram[21312]  = 1;
  ram[21313]  = 1;
  ram[21314]  = 1;
  ram[21315]  = 1;
  ram[21316]  = 1;
  ram[21317]  = 1;
  ram[21318]  = 1;
  ram[21319]  = 1;
  ram[21320]  = 1;
  ram[21321]  = 1;
  ram[21322]  = 1;
  ram[21323]  = 1;
  ram[21324]  = 1;
  ram[21325]  = 1;
  ram[21326]  = 1;
  ram[21327]  = 1;
  ram[21328]  = 1;
  ram[21329]  = 1;
  ram[21330]  = 1;
  ram[21331]  = 1;
  ram[21332]  = 1;
  ram[21333]  = 1;
  ram[21334]  = 1;
  ram[21335]  = 1;
  ram[21336]  = 1;
  ram[21337]  = 1;
  ram[21338]  = 1;
  ram[21339]  = 1;
  ram[21340]  = 1;
  ram[21341]  = 1;
  ram[21342]  = 1;
  ram[21343]  = 1;
  ram[21344]  = 1;
  ram[21345]  = 0;
  ram[21346]  = 1;
  ram[21347]  = 1;
  ram[21348]  = 1;
  ram[21349]  = 1;
  ram[21350]  = 0;
  ram[21351]  = 0;
  ram[21352]  = 1;
  ram[21353]  = 1;
  ram[21354]  = 1;
  ram[21355]  = 0;
  ram[21356]  = 1;
  ram[21357]  = 1;
  ram[21358]  = 1;
  ram[21359]  = 1;
  ram[21360]  = 1;
  ram[21361]  = 0;
  ram[21362]  = 1;
  ram[21363]  = 1;
  ram[21364]  = 1;
  ram[21365]  = 1;
  ram[21366]  = 1;
  ram[21367]  = 0;
  ram[21368]  = 1;
  ram[21369]  = 1;
  ram[21370]  = 0;
  ram[21371]  = 1;
  ram[21372]  = 1;
  ram[21373]  = 1;
  ram[21374]  = 1;
  ram[21375]  = 1;
  ram[21376]  = 1;
  ram[21377]  = 0;
  ram[21378]  = 0;
  ram[21379]  = 1;
  ram[21380]  = 1;
  ram[21381]  = 1;
  ram[21382]  = 1;
  ram[21383]  = 1;
  ram[21384]  = 1;
  ram[21385]  = 1;
  ram[21386]  = 1;
  ram[21387]  = 1;
  ram[21388]  = 1;
  ram[21389]  = 1;
  ram[21390]  = 1;
  ram[21391]  = 0;
  ram[21392]  = 1;
  ram[21393]  = 1;
  ram[21394]  = 1;
  ram[21395]  = 1;
  ram[21396]  = 1;
  ram[21397]  = 0;
  ram[21398]  = 1;
  ram[21399]  = 1;
  ram[21400]  = 1;
  ram[21401]  = 1;
  ram[21402]  = 1;
  ram[21403]  = 0;
  ram[21404]  = 1;
  ram[21405]  = 1;
  ram[21406]  = 1;
  ram[21407]  = 0;
  ram[21408]  = 1;
  ram[21409]  = 1;
  ram[21410]  = 1;
  ram[21411]  = 1;
  ram[21412]  = 1;
  ram[21413]  = 0;
  ram[21414]  = 1;
  ram[21415]  = 1;
  ram[21416]  = 1;
  ram[21417]  = 1;
  ram[21418]  = 1;
  ram[21419]  = 1;
  ram[21420]  = 1;
  ram[21421]  = 1;
  ram[21422]  = 0;
  ram[21423]  = 0;
  ram[21424]  = 0;
  ram[21425]  = 0;
  ram[21426]  = 0;
  ram[21427]  = 1;
  ram[21428]  = 1;
  ram[21429]  = 1;
  ram[21430]  = 1;
  ram[21431]  = 1;
  ram[21432]  = 0;
  ram[21433]  = 1;
  ram[21434]  = 1;
  ram[21435]  = 1;
  ram[21436]  = 1;
  ram[21437]  = 1;
  ram[21438]  = 0;
  ram[21439]  = 1;
  ram[21440]  = 1;
  ram[21441]  = 1;
  ram[21442]  = 0;
  ram[21443]  = 0;
  ram[21444]  = 1;
  ram[21445]  = 1;
  ram[21446]  = 1;
  ram[21447]  = 1;
  ram[21448]  = 0;
  ram[21449]  = 1;
  ram[21450]  = 1;
  ram[21451]  = 1;
  ram[21452]  = 1;
  ram[21453]  = 1;
  ram[21454]  = 0;
  ram[21455]  = 1;
  ram[21456]  = 1;
  ram[21457]  = 1;
  ram[21458]  = 1;
  ram[21459]  = 1;
  ram[21460]  = 1;
  ram[21461]  = 0;
  ram[21462]  = 1;
  ram[21463]  = 1;
  ram[21464]  = 1;
  ram[21465]  = 0;
  ram[21466]  = 1;
  ram[21467]  = 1;
  ram[21468]  = 1;
  ram[21469]  = 1;
  ram[21470]  = 1;
  ram[21471]  = 0;
  ram[21472]  = 1;
  ram[21473]  = 1;
  ram[21474]  = 1;
  ram[21475]  = 1;
  ram[21476]  = 1;
  ram[21477]  = 1;
  ram[21478]  = 1;
  ram[21479]  = 1;
  ram[21480]  = 0;
  ram[21481]  = 1;
  ram[21482]  = 1;
  ram[21483]  = 1;
  ram[21484]  = 1;
  ram[21485]  = 0;
  ram[21486]  = 0;
  ram[21487]  = 1;
  ram[21488]  = 1;
  ram[21489]  = 1;
  ram[21490]  = 1;
  ram[21491]  = 1;
  ram[21492]  = 0;
  ram[21493]  = 0;
  ram[21494]  = 1;
  ram[21495]  = 1;
  ram[21496]  = 1;
  ram[21497]  = 1;
  ram[21498]  = 1;
  ram[21499]  = 1;
  ram[21500]  = 1;
  ram[21501]  = 0;
  ram[21502]  = 0;
  ram[21503]  = 1;
  ram[21504]  = 1;
  ram[21505]  = 1;
  ram[21506]  = 1;
  ram[21507]  = 0;
  ram[21508]  = 1;
  ram[21509]  = 1;
  ram[21510]  = 1;
  ram[21511]  = 1;
  ram[21512]  = 1;
  ram[21513]  = 1;
  ram[21514]  = 0;
  ram[21515]  = 1;
  ram[21516]  = 0;
  ram[21517]  = 0;
  ram[21518]  = 1;
  ram[21519]  = 1;
  ram[21520]  = 1;
  ram[21521]  = 1;
  ram[21522]  = 1;
  ram[21523]  = 1;
  ram[21524]  = 1;
  ram[21525]  = 0;
  ram[21526]  = 1;
  ram[21527]  = 1;
  ram[21528]  = 1;
  ram[21529]  = 1;
  ram[21530]  = 1;
  ram[21531]  = 1;
  ram[21532]  = 1;
  ram[21533]  = 1;
  ram[21534]  = 1;
  ram[21535]  = 1;
  ram[21536]  = 0;
  ram[21537]  = 1;
  ram[21538]  = 1;
  ram[21539]  = 1;
  ram[21540]  = 0;
  ram[21541]  = 1;
  ram[21542]  = 1;
  ram[21543]  = 1;
  ram[21544]  = 1;
  ram[21545]  = 1;
  ram[21546]  = 0;
  ram[21547]  = 0;
  ram[21548]  = 1;
  ram[21549]  = 1;
  ram[21550]  = 1;
  ram[21551]  = 1;
  ram[21552]  = 1;
  ram[21553]  = 1;
  ram[21554]  = 1;
  ram[21555]  = 1;
  ram[21556]  = 1;
  ram[21557]  = 1;
  ram[21558]  = 1;
  ram[21559]  = 1;
  ram[21560]  = 1;
  ram[21561]  = 1;
  ram[21562]  = 1;
  ram[21563]  = 1;
  ram[21564]  = 1;
  ram[21565]  = 1;
  ram[21566]  = 1;
  ram[21567]  = 1;
  ram[21568]  = 1;
  ram[21569]  = 1;
  ram[21570]  = 1;
  ram[21571]  = 1;
  ram[21572]  = 1;
  ram[21573]  = 1;
  ram[21574]  = 1;
  ram[21575]  = 1;
  ram[21576]  = 1;
  ram[21577]  = 1;
  ram[21578]  = 1;
  ram[21579]  = 1;
  ram[21580]  = 1;
  ram[21581]  = 1;
  ram[21582]  = 1;
  ram[21583]  = 1;
  ram[21584]  = 1;
  ram[21585]  = 1;
  ram[21586]  = 1;
  ram[21587]  = 1;
  ram[21588]  = 1;
  ram[21589]  = 1;
  ram[21590]  = 1;
  ram[21591]  = 1;
  ram[21592]  = 1;
  ram[21593]  = 1;
  ram[21594]  = 1;
  ram[21595]  = 1;
  ram[21596]  = 1;
  ram[21597]  = 1;
  ram[21598]  = 1;
  ram[21599]  = 1;
  ram[21600]  = 1;
  ram[21601]  = 1;
  ram[21602]  = 1;
  ram[21603]  = 1;
  ram[21604]  = 1;
  ram[21605]  = 1;
  ram[21606]  = 1;
  ram[21607]  = 1;
  ram[21608]  = 1;
  ram[21609]  = 1;
  ram[21610]  = 1;
  ram[21611]  = 1;
  ram[21612]  = 1;
  ram[21613]  = 1;
  ram[21614]  = 1;
  ram[21615]  = 1;
  ram[21616]  = 1;
  ram[21617]  = 1;
  ram[21618]  = 1;
  ram[21619]  = 1;
  ram[21620]  = 1;
  ram[21621]  = 1;
  ram[21622]  = 1;
  ram[21623]  = 1;
  ram[21624]  = 1;
  ram[21625]  = 1;
  ram[21626]  = 1;
  ram[21627]  = 1;
  ram[21628]  = 1;
  ram[21629]  = 1;
  ram[21630]  = 1;
  ram[21631]  = 1;
  ram[21632]  = 1;
  ram[21633]  = 1;
  ram[21634]  = 1;
  ram[21635]  = 1;
  ram[21636]  = 1;
  ram[21637]  = 1;
  ram[21638]  = 1;
  ram[21639]  = 1;
  ram[21640]  = 1;
  ram[21641]  = 1;
  ram[21642]  = 1;
  ram[21643]  = 1;
  ram[21644]  = 1;
  ram[21645]  = 0;
  ram[21646]  = 1;
  ram[21647]  = 1;
  ram[21648]  = 1;
  ram[21649]  = 0;
  ram[21650]  = 0;
  ram[21651]  = 1;
  ram[21652]  = 1;
  ram[21653]  = 1;
  ram[21654]  = 1;
  ram[21655]  = 0;
  ram[21656]  = 1;
  ram[21657]  = 1;
  ram[21658]  = 1;
  ram[21659]  = 1;
  ram[21660]  = 1;
  ram[21661]  = 0;
  ram[21662]  = 1;
  ram[21663]  = 1;
  ram[21664]  = 1;
  ram[21665]  = 1;
  ram[21666]  = 1;
  ram[21667]  = 0;
  ram[21668]  = 1;
  ram[21669]  = 1;
  ram[21670]  = 0;
  ram[21671]  = 1;
  ram[21672]  = 1;
  ram[21673]  = 1;
  ram[21674]  = 1;
  ram[21675]  = 1;
  ram[21676]  = 1;
  ram[21677]  = 1;
  ram[21678]  = 0;
  ram[21679]  = 1;
  ram[21680]  = 1;
  ram[21681]  = 1;
  ram[21682]  = 1;
  ram[21683]  = 1;
  ram[21684]  = 1;
  ram[21685]  = 1;
  ram[21686]  = 1;
  ram[21687]  = 1;
  ram[21688]  = 1;
  ram[21689]  = 1;
  ram[21690]  = 1;
  ram[21691]  = 0;
  ram[21692]  = 1;
  ram[21693]  = 1;
  ram[21694]  = 1;
  ram[21695]  = 1;
  ram[21696]  = 1;
  ram[21697]  = 0;
  ram[21698]  = 1;
  ram[21699]  = 1;
  ram[21700]  = 1;
  ram[21701]  = 1;
  ram[21702]  = 1;
  ram[21703]  = 0;
  ram[21704]  = 1;
  ram[21705]  = 1;
  ram[21706]  = 0;
  ram[21707]  = 0;
  ram[21708]  = 1;
  ram[21709]  = 1;
  ram[21710]  = 1;
  ram[21711]  = 1;
  ram[21712]  = 1;
  ram[21713]  = 0;
  ram[21714]  = 1;
  ram[21715]  = 1;
  ram[21716]  = 1;
  ram[21717]  = 1;
  ram[21718]  = 1;
  ram[21719]  = 1;
  ram[21720]  = 1;
  ram[21721]  = 1;
  ram[21722]  = 0;
  ram[21723]  = 1;
  ram[21724]  = 1;
  ram[21725]  = 1;
  ram[21726]  = 0;
  ram[21727]  = 0;
  ram[21728]  = 1;
  ram[21729]  = 1;
  ram[21730]  = 1;
  ram[21731]  = 1;
  ram[21732]  = 0;
  ram[21733]  = 1;
  ram[21734]  = 1;
  ram[21735]  = 1;
  ram[21736]  = 1;
  ram[21737]  = 1;
  ram[21738]  = 0;
  ram[21739]  = 1;
  ram[21740]  = 1;
  ram[21741]  = 1;
  ram[21742]  = 0;
  ram[21743]  = 0;
  ram[21744]  = 1;
  ram[21745]  = 1;
  ram[21746]  = 1;
  ram[21747]  = 1;
  ram[21748]  = 0;
  ram[21749]  = 1;
  ram[21750]  = 1;
  ram[21751]  = 1;
  ram[21752]  = 1;
  ram[21753]  = 0;
  ram[21754]  = 0;
  ram[21755]  = 1;
  ram[21756]  = 1;
  ram[21757]  = 1;
  ram[21758]  = 1;
  ram[21759]  = 1;
  ram[21760]  = 1;
  ram[21761]  = 0;
  ram[21762]  = 1;
  ram[21763]  = 1;
  ram[21764]  = 0;
  ram[21765]  = 0;
  ram[21766]  = 1;
  ram[21767]  = 1;
  ram[21768]  = 1;
  ram[21769]  = 1;
  ram[21770]  = 1;
  ram[21771]  = 0;
  ram[21772]  = 1;
  ram[21773]  = 1;
  ram[21774]  = 1;
  ram[21775]  = 1;
  ram[21776]  = 1;
  ram[21777]  = 1;
  ram[21778]  = 1;
  ram[21779]  = 1;
  ram[21780]  = 0;
  ram[21781]  = 1;
  ram[21782]  = 1;
  ram[21783]  = 1;
  ram[21784]  = 1;
  ram[21785]  = 0;
  ram[21786]  = 1;
  ram[21787]  = 1;
  ram[21788]  = 1;
  ram[21789]  = 1;
  ram[21790]  = 1;
  ram[21791]  = 1;
  ram[21792]  = 1;
  ram[21793]  = 0;
  ram[21794]  = 1;
  ram[21795]  = 1;
  ram[21796]  = 1;
  ram[21797]  = 1;
  ram[21798]  = 1;
  ram[21799]  = 1;
  ram[21800]  = 1;
  ram[21801]  = 0;
  ram[21802]  = 0;
  ram[21803]  = 1;
  ram[21804]  = 1;
  ram[21805]  = 1;
  ram[21806]  = 1;
  ram[21807]  = 0;
  ram[21808]  = 1;
  ram[21809]  = 1;
  ram[21810]  = 1;
  ram[21811]  = 1;
  ram[21812]  = 1;
  ram[21813]  = 1;
  ram[21814]  = 0;
  ram[21815]  = 1;
  ram[21816]  = 1;
  ram[21817]  = 0;
  ram[21818]  = 1;
  ram[21819]  = 1;
  ram[21820]  = 1;
  ram[21821]  = 1;
  ram[21822]  = 1;
  ram[21823]  = 1;
  ram[21824]  = 1;
  ram[21825]  = 0;
  ram[21826]  = 1;
  ram[21827]  = 1;
  ram[21828]  = 1;
  ram[21829]  = 1;
  ram[21830]  = 1;
  ram[21831]  = 1;
  ram[21832]  = 1;
  ram[21833]  = 1;
  ram[21834]  = 1;
  ram[21835]  = 1;
  ram[21836]  = 0;
  ram[21837]  = 1;
  ram[21838]  = 1;
  ram[21839]  = 1;
  ram[21840]  = 0;
  ram[21841]  = 1;
  ram[21842]  = 1;
  ram[21843]  = 1;
  ram[21844]  = 1;
  ram[21845]  = 1;
  ram[21846]  = 0;
  ram[21847]  = 0;
  ram[21848]  = 1;
  ram[21849]  = 1;
  ram[21850]  = 1;
  ram[21851]  = 1;
  ram[21852]  = 1;
  ram[21853]  = 1;
  ram[21854]  = 1;
  ram[21855]  = 1;
  ram[21856]  = 1;
  ram[21857]  = 1;
  ram[21858]  = 1;
  ram[21859]  = 1;
  ram[21860]  = 1;
  ram[21861]  = 1;
  ram[21862]  = 1;
  ram[21863]  = 1;
  ram[21864]  = 1;
  ram[21865]  = 1;
  ram[21866]  = 1;
  ram[21867]  = 1;
  ram[21868]  = 1;
  ram[21869]  = 1;
  ram[21870]  = 1;
  ram[21871]  = 1;
  ram[21872]  = 1;
  ram[21873]  = 1;
  ram[21874]  = 1;
  ram[21875]  = 1;
  ram[21876]  = 1;
  ram[21877]  = 1;
  ram[21878]  = 1;
  ram[21879]  = 1;
  ram[21880]  = 1;
  ram[21881]  = 1;
  ram[21882]  = 1;
  ram[21883]  = 1;
  ram[21884]  = 1;
  ram[21885]  = 1;
  ram[21886]  = 1;
  ram[21887]  = 1;
  ram[21888]  = 1;
  ram[21889]  = 1;
  ram[21890]  = 1;
  ram[21891]  = 1;
  ram[21892]  = 1;
  ram[21893]  = 1;
  ram[21894]  = 1;
  ram[21895]  = 1;
  ram[21896]  = 1;
  ram[21897]  = 1;
  ram[21898]  = 1;
  ram[21899]  = 1;
  ram[21900]  = 1;
  ram[21901]  = 1;
  ram[21902]  = 1;
  ram[21903]  = 1;
  ram[21904]  = 1;
  ram[21905]  = 1;
  ram[21906]  = 1;
  ram[21907]  = 1;
  ram[21908]  = 1;
  ram[21909]  = 1;
  ram[21910]  = 1;
  ram[21911]  = 1;
  ram[21912]  = 1;
  ram[21913]  = 1;
  ram[21914]  = 1;
  ram[21915]  = 1;
  ram[21916]  = 1;
  ram[21917]  = 1;
  ram[21918]  = 1;
  ram[21919]  = 1;
  ram[21920]  = 1;
  ram[21921]  = 1;
  ram[21922]  = 1;
  ram[21923]  = 1;
  ram[21924]  = 1;
  ram[21925]  = 1;
  ram[21926]  = 1;
  ram[21927]  = 1;
  ram[21928]  = 1;
  ram[21929]  = 1;
  ram[21930]  = 1;
  ram[21931]  = 1;
  ram[21932]  = 1;
  ram[21933]  = 1;
  ram[21934]  = 1;
  ram[21935]  = 1;
  ram[21936]  = 1;
  ram[21937]  = 1;
  ram[21938]  = 1;
  ram[21939]  = 1;
  ram[21940]  = 1;
  ram[21941]  = 1;
  ram[21942]  = 1;
  ram[21943]  = 1;
  ram[21944]  = 1;
  ram[21945]  = 0;
  ram[21946]  = 0;
  ram[21947]  = 0;
  ram[21948]  = 0;
  ram[21949]  = 0;
  ram[21950]  = 0;
  ram[21951]  = 1;
  ram[21952]  = 1;
  ram[21953]  = 1;
  ram[21954]  = 1;
  ram[21955]  = 0;
  ram[21956]  = 1;
  ram[21957]  = 1;
  ram[21958]  = 1;
  ram[21959]  = 1;
  ram[21960]  = 1;
  ram[21961]  = 0;
  ram[21962]  = 1;
  ram[21963]  = 1;
  ram[21964]  = 1;
  ram[21965]  = 1;
  ram[21966]  = 1;
  ram[21967]  = 0;
  ram[21968]  = 1;
  ram[21969]  = 1;
  ram[21970]  = 0;
  ram[21971]  = 0;
  ram[21972]  = 1;
  ram[21973]  = 1;
  ram[21974]  = 1;
  ram[21975]  = 1;
  ram[21976]  = 1;
  ram[21977]  = 1;
  ram[21978]  = 0;
  ram[21979]  = 0;
  ram[21980]  = 1;
  ram[21981]  = 1;
  ram[21982]  = 1;
  ram[21983]  = 1;
  ram[21984]  = 1;
  ram[21985]  = 1;
  ram[21986]  = 1;
  ram[21987]  = 1;
  ram[21988]  = 1;
  ram[21989]  = 1;
  ram[21990]  = 1;
  ram[21991]  = 0;
  ram[21992]  = 1;
  ram[21993]  = 1;
  ram[21994]  = 1;
  ram[21995]  = 1;
  ram[21996]  = 1;
  ram[21997]  = 0;
  ram[21998]  = 1;
  ram[21999]  = 1;
  ram[22000]  = 1;
  ram[22001]  = 1;
  ram[22002]  = 1;
  ram[22003]  = 0;
  ram[22004]  = 1;
  ram[22005]  = 1;
  ram[22006]  = 0;
  ram[22007]  = 0;
  ram[22008]  = 1;
  ram[22009]  = 1;
  ram[22010]  = 1;
  ram[22011]  = 1;
  ram[22012]  = 1;
  ram[22013]  = 0;
  ram[22014]  = 1;
  ram[22015]  = 1;
  ram[22016]  = 1;
  ram[22017]  = 1;
  ram[22018]  = 1;
  ram[22019]  = 1;
  ram[22020]  = 1;
  ram[22021]  = 1;
  ram[22022]  = 0;
  ram[22023]  = 1;
  ram[22024]  = 1;
  ram[22025]  = 1;
  ram[22026]  = 1;
  ram[22027]  = 1;
  ram[22028]  = 0;
  ram[22029]  = 1;
  ram[22030]  = 1;
  ram[22031]  = 1;
  ram[22032]  = 0;
  ram[22033]  = 1;
  ram[22034]  = 1;
  ram[22035]  = 1;
  ram[22036]  = 1;
  ram[22037]  = 1;
  ram[22038]  = 0;
  ram[22039]  = 1;
  ram[22040]  = 1;
  ram[22041]  = 1;
  ram[22042]  = 0;
  ram[22043]  = 0;
  ram[22044]  = 1;
  ram[22045]  = 1;
  ram[22046]  = 1;
  ram[22047]  = 1;
  ram[22048]  = 0;
  ram[22049]  = 1;
  ram[22050]  = 1;
  ram[22051]  = 1;
  ram[22052]  = 1;
  ram[22053]  = 0;
  ram[22054]  = 0;
  ram[22055]  = 1;
  ram[22056]  = 1;
  ram[22057]  = 1;
  ram[22058]  = 1;
  ram[22059]  = 1;
  ram[22060]  = 1;
  ram[22061]  = 0;
  ram[22062]  = 1;
  ram[22063]  = 1;
  ram[22064]  = 0;
  ram[22065]  = 0;
  ram[22066]  = 1;
  ram[22067]  = 1;
  ram[22068]  = 1;
  ram[22069]  = 1;
  ram[22070]  = 1;
  ram[22071]  = 0;
  ram[22072]  = 1;
  ram[22073]  = 1;
  ram[22074]  = 1;
  ram[22075]  = 1;
  ram[22076]  = 1;
  ram[22077]  = 1;
  ram[22078]  = 1;
  ram[22079]  = 1;
  ram[22080]  = 0;
  ram[22081]  = 1;
  ram[22082]  = 1;
  ram[22083]  = 1;
  ram[22084]  = 1;
  ram[22085]  = 0;
  ram[22086]  = 1;
  ram[22087]  = 1;
  ram[22088]  = 1;
  ram[22089]  = 1;
  ram[22090]  = 1;
  ram[22091]  = 1;
  ram[22092]  = 1;
  ram[22093]  = 0;
  ram[22094]  = 1;
  ram[22095]  = 1;
  ram[22096]  = 1;
  ram[22097]  = 1;
  ram[22098]  = 1;
  ram[22099]  = 1;
  ram[22100]  = 1;
  ram[22101]  = 0;
  ram[22102]  = 0;
  ram[22103]  = 1;
  ram[22104]  = 1;
  ram[22105]  = 1;
  ram[22106]  = 1;
  ram[22107]  = 0;
  ram[22108]  = 1;
  ram[22109]  = 1;
  ram[22110]  = 1;
  ram[22111]  = 1;
  ram[22112]  = 1;
  ram[22113]  = 1;
  ram[22114]  = 0;
  ram[22115]  = 1;
  ram[22116]  = 1;
  ram[22117]  = 0;
  ram[22118]  = 0;
  ram[22119]  = 1;
  ram[22120]  = 1;
  ram[22121]  = 1;
  ram[22122]  = 1;
  ram[22123]  = 1;
  ram[22124]  = 1;
  ram[22125]  = 0;
  ram[22126]  = 1;
  ram[22127]  = 1;
  ram[22128]  = 1;
  ram[22129]  = 1;
  ram[22130]  = 1;
  ram[22131]  = 1;
  ram[22132]  = 1;
  ram[22133]  = 0;
  ram[22134]  = 0;
  ram[22135]  = 0;
  ram[22136]  = 0;
  ram[22137]  = 1;
  ram[22138]  = 1;
  ram[22139]  = 1;
  ram[22140]  = 0;
  ram[22141]  = 1;
  ram[22142]  = 1;
  ram[22143]  = 1;
  ram[22144]  = 1;
  ram[22145]  = 1;
  ram[22146]  = 0;
  ram[22147]  = 0;
  ram[22148]  = 1;
  ram[22149]  = 1;
  ram[22150]  = 1;
  ram[22151]  = 1;
  ram[22152]  = 1;
  ram[22153]  = 1;
  ram[22154]  = 1;
  ram[22155]  = 1;
  ram[22156]  = 1;
  ram[22157]  = 1;
  ram[22158]  = 1;
  ram[22159]  = 1;
  ram[22160]  = 1;
  ram[22161]  = 1;
  ram[22162]  = 1;
  ram[22163]  = 1;
  ram[22164]  = 1;
  ram[22165]  = 1;
  ram[22166]  = 1;
  ram[22167]  = 1;
  ram[22168]  = 1;
  ram[22169]  = 1;
  ram[22170]  = 1;
  ram[22171]  = 1;
  ram[22172]  = 1;
  ram[22173]  = 1;
  ram[22174]  = 1;
  ram[22175]  = 1;
  ram[22176]  = 1;
  ram[22177]  = 1;
  ram[22178]  = 1;
  ram[22179]  = 1;
  ram[22180]  = 1;
  ram[22181]  = 1;
  ram[22182]  = 1;
  ram[22183]  = 1;
  ram[22184]  = 1;
  ram[22185]  = 1;
  ram[22186]  = 1;
  ram[22187]  = 1;
  ram[22188]  = 1;
  ram[22189]  = 1;
  ram[22190]  = 1;
  ram[22191]  = 1;
  ram[22192]  = 1;
  ram[22193]  = 1;
  ram[22194]  = 1;
  ram[22195]  = 1;
  ram[22196]  = 1;
  ram[22197]  = 1;
  ram[22198]  = 1;
  ram[22199]  = 1;
  ram[22200]  = 1;
  ram[22201]  = 1;
  ram[22202]  = 1;
  ram[22203]  = 1;
  ram[22204]  = 1;
  ram[22205]  = 1;
  ram[22206]  = 1;
  ram[22207]  = 1;
  ram[22208]  = 1;
  ram[22209]  = 1;
  ram[22210]  = 1;
  ram[22211]  = 1;
  ram[22212]  = 1;
  ram[22213]  = 1;
  ram[22214]  = 1;
  ram[22215]  = 1;
  ram[22216]  = 1;
  ram[22217]  = 1;
  ram[22218]  = 1;
  ram[22219]  = 1;
  ram[22220]  = 1;
  ram[22221]  = 1;
  ram[22222]  = 1;
  ram[22223]  = 1;
  ram[22224]  = 1;
  ram[22225]  = 1;
  ram[22226]  = 1;
  ram[22227]  = 1;
  ram[22228]  = 1;
  ram[22229]  = 1;
  ram[22230]  = 1;
  ram[22231]  = 1;
  ram[22232]  = 1;
  ram[22233]  = 1;
  ram[22234]  = 1;
  ram[22235]  = 1;
  ram[22236]  = 1;
  ram[22237]  = 1;
  ram[22238]  = 1;
  ram[22239]  = 1;
  ram[22240]  = 1;
  ram[22241]  = 1;
  ram[22242]  = 1;
  ram[22243]  = 1;
  ram[22244]  = 1;
  ram[22245]  = 0;
  ram[22246]  = 1;
  ram[22247]  = 1;
  ram[22248]  = 1;
  ram[22249]  = 1;
  ram[22250]  = 1;
  ram[22251]  = 1;
  ram[22252]  = 1;
  ram[22253]  = 1;
  ram[22254]  = 1;
  ram[22255]  = 0;
  ram[22256]  = 1;
  ram[22257]  = 1;
  ram[22258]  = 1;
  ram[22259]  = 1;
  ram[22260]  = 1;
  ram[22261]  = 0;
  ram[22262]  = 0;
  ram[22263]  = 0;
  ram[22264]  = 0;
  ram[22265]  = 0;
  ram[22266]  = 0;
  ram[22267]  = 0;
  ram[22268]  = 0;
  ram[22269]  = 1;
  ram[22270]  = 1;
  ram[22271]  = 0;
  ram[22272]  = 0;
  ram[22273]  = 0;
  ram[22274]  = 1;
  ram[22275]  = 1;
  ram[22276]  = 1;
  ram[22277]  = 1;
  ram[22278]  = 1;
  ram[22279]  = 0;
  ram[22280]  = 0;
  ram[22281]  = 0;
  ram[22282]  = 1;
  ram[22283]  = 1;
  ram[22284]  = 1;
  ram[22285]  = 1;
  ram[22286]  = 1;
  ram[22287]  = 1;
  ram[22288]  = 1;
  ram[22289]  = 1;
  ram[22290]  = 1;
  ram[22291]  = 0;
  ram[22292]  = 1;
  ram[22293]  = 1;
  ram[22294]  = 1;
  ram[22295]  = 1;
  ram[22296]  = 1;
  ram[22297]  = 0;
  ram[22298]  = 1;
  ram[22299]  = 1;
  ram[22300]  = 1;
  ram[22301]  = 1;
  ram[22302]  = 1;
  ram[22303]  = 0;
  ram[22304]  = 1;
  ram[22305]  = 1;
  ram[22306]  = 0;
  ram[22307]  = 0;
  ram[22308]  = 0;
  ram[22309]  = 0;
  ram[22310]  = 0;
  ram[22311]  = 0;
  ram[22312]  = 0;
  ram[22313]  = 0;
  ram[22314]  = 1;
  ram[22315]  = 1;
  ram[22316]  = 1;
  ram[22317]  = 1;
  ram[22318]  = 1;
  ram[22319]  = 1;
  ram[22320]  = 1;
  ram[22321]  = 1;
  ram[22322]  = 0;
  ram[22323]  = 1;
  ram[22324]  = 1;
  ram[22325]  = 1;
  ram[22326]  = 1;
  ram[22327]  = 1;
  ram[22328]  = 0;
  ram[22329]  = 1;
  ram[22330]  = 1;
  ram[22331]  = 1;
  ram[22332]  = 0;
  ram[22333]  = 1;
  ram[22334]  = 1;
  ram[22335]  = 1;
  ram[22336]  = 1;
  ram[22337]  = 1;
  ram[22338]  = 0;
  ram[22339]  = 1;
  ram[22340]  = 1;
  ram[22341]  = 1;
  ram[22342]  = 0;
  ram[22343]  = 0;
  ram[22344]  = 1;
  ram[22345]  = 1;
  ram[22346]  = 1;
  ram[22347]  = 1;
  ram[22348]  = 0;
  ram[22349]  = 1;
  ram[22350]  = 1;
  ram[22351]  = 1;
  ram[22352]  = 1;
  ram[22353]  = 0;
  ram[22354]  = 0;
  ram[22355]  = 1;
  ram[22356]  = 1;
  ram[22357]  = 1;
  ram[22358]  = 1;
  ram[22359]  = 1;
  ram[22360]  = 1;
  ram[22361]  = 0;
  ram[22362]  = 1;
  ram[22363]  = 1;
  ram[22364]  = 0;
  ram[22365]  = 0;
  ram[22366]  = 1;
  ram[22367]  = 1;
  ram[22368]  = 1;
  ram[22369]  = 1;
  ram[22370]  = 1;
  ram[22371]  = 0;
  ram[22372]  = 1;
  ram[22373]  = 1;
  ram[22374]  = 1;
  ram[22375]  = 1;
  ram[22376]  = 1;
  ram[22377]  = 1;
  ram[22378]  = 1;
  ram[22379]  = 1;
  ram[22380]  = 0;
  ram[22381]  = 1;
  ram[22382]  = 1;
  ram[22383]  = 1;
  ram[22384]  = 1;
  ram[22385]  = 0;
  ram[22386]  = 1;
  ram[22387]  = 1;
  ram[22388]  = 1;
  ram[22389]  = 1;
  ram[22390]  = 1;
  ram[22391]  = 1;
  ram[22392]  = 1;
  ram[22393]  = 0;
  ram[22394]  = 1;
  ram[22395]  = 1;
  ram[22396]  = 1;
  ram[22397]  = 1;
  ram[22398]  = 1;
  ram[22399]  = 1;
  ram[22400]  = 1;
  ram[22401]  = 0;
  ram[22402]  = 0;
  ram[22403]  = 1;
  ram[22404]  = 1;
  ram[22405]  = 1;
  ram[22406]  = 1;
  ram[22407]  = 0;
  ram[22408]  = 0;
  ram[22409]  = 0;
  ram[22410]  = 0;
  ram[22411]  = 0;
  ram[22412]  = 0;
  ram[22413]  = 0;
  ram[22414]  = 0;
  ram[22415]  = 1;
  ram[22416]  = 1;
  ram[22417]  = 1;
  ram[22418]  = 0;
  ram[22419]  = 0;
  ram[22420]  = 0;
  ram[22421]  = 1;
  ram[22422]  = 1;
  ram[22423]  = 1;
  ram[22424]  = 1;
  ram[22425]  = 0;
  ram[22426]  = 1;
  ram[22427]  = 1;
  ram[22428]  = 1;
  ram[22429]  = 1;
  ram[22430]  = 1;
  ram[22431]  = 0;
  ram[22432]  = 0;
  ram[22433]  = 0;
  ram[22434]  = 0;
  ram[22435]  = 0;
  ram[22436]  = 0;
  ram[22437]  = 1;
  ram[22438]  = 1;
  ram[22439]  = 1;
  ram[22440]  = 0;
  ram[22441]  = 1;
  ram[22442]  = 1;
  ram[22443]  = 1;
  ram[22444]  = 1;
  ram[22445]  = 1;
  ram[22446]  = 0;
  ram[22447]  = 0;
  ram[22448]  = 1;
  ram[22449]  = 1;
  ram[22450]  = 1;
  ram[22451]  = 1;
  ram[22452]  = 1;
  ram[22453]  = 1;
  ram[22454]  = 1;
  ram[22455]  = 1;
  ram[22456]  = 1;
  ram[22457]  = 1;
  ram[22458]  = 1;
  ram[22459]  = 1;
  ram[22460]  = 1;
  ram[22461]  = 1;
  ram[22462]  = 1;
  ram[22463]  = 1;
  ram[22464]  = 1;
  ram[22465]  = 1;
  ram[22466]  = 1;
  ram[22467]  = 1;
  ram[22468]  = 1;
  ram[22469]  = 1;
  ram[22470]  = 1;
  ram[22471]  = 1;
  ram[22472]  = 1;
  ram[22473]  = 1;
  ram[22474]  = 1;
  ram[22475]  = 1;
  ram[22476]  = 1;
  ram[22477]  = 1;
  ram[22478]  = 1;
  ram[22479]  = 1;
  ram[22480]  = 1;
  ram[22481]  = 1;
  ram[22482]  = 1;
  ram[22483]  = 1;
  ram[22484]  = 1;
  ram[22485]  = 1;
  ram[22486]  = 1;
  ram[22487]  = 1;
  ram[22488]  = 1;
  ram[22489]  = 1;
  ram[22490]  = 1;
  ram[22491]  = 1;
  ram[22492]  = 1;
  ram[22493]  = 1;
  ram[22494]  = 1;
  ram[22495]  = 1;
  ram[22496]  = 1;
  ram[22497]  = 1;
  ram[22498]  = 1;
  ram[22499]  = 1;
  ram[22500]  = 1;
  ram[22501]  = 1;
  ram[22502]  = 1;
  ram[22503]  = 1;
  ram[22504]  = 1;
  ram[22505]  = 1;
  ram[22506]  = 1;
  ram[22507]  = 1;
  ram[22508]  = 1;
  ram[22509]  = 1;
  ram[22510]  = 1;
  ram[22511]  = 1;
  ram[22512]  = 1;
  ram[22513]  = 1;
  ram[22514]  = 1;
  ram[22515]  = 1;
  ram[22516]  = 1;
  ram[22517]  = 1;
  ram[22518]  = 1;
  ram[22519]  = 1;
  ram[22520]  = 1;
  ram[22521]  = 1;
  ram[22522]  = 1;
  ram[22523]  = 1;
  ram[22524]  = 1;
  ram[22525]  = 1;
  ram[22526]  = 1;
  ram[22527]  = 1;
  ram[22528]  = 1;
  ram[22529]  = 1;
  ram[22530]  = 1;
  ram[22531]  = 1;
  ram[22532]  = 1;
  ram[22533]  = 1;
  ram[22534]  = 1;
  ram[22535]  = 1;
  ram[22536]  = 1;
  ram[22537]  = 1;
  ram[22538]  = 1;
  ram[22539]  = 1;
  ram[22540]  = 1;
  ram[22541]  = 1;
  ram[22542]  = 1;
  ram[22543]  = 1;
  ram[22544]  = 1;
  ram[22545]  = 0;
  ram[22546]  = 1;
  ram[22547]  = 1;
  ram[22548]  = 1;
  ram[22549]  = 1;
  ram[22550]  = 1;
  ram[22551]  = 1;
  ram[22552]  = 1;
  ram[22553]  = 1;
  ram[22554]  = 1;
  ram[22555]  = 0;
  ram[22556]  = 1;
  ram[22557]  = 1;
  ram[22558]  = 1;
  ram[22559]  = 1;
  ram[22560]  = 1;
  ram[22561]  = 0;
  ram[22562]  = 1;
  ram[22563]  = 1;
  ram[22564]  = 1;
  ram[22565]  = 1;
  ram[22566]  = 1;
  ram[22567]  = 1;
  ram[22568]  = 1;
  ram[22569]  = 1;
  ram[22570]  = 1;
  ram[22571]  = 1;
  ram[22572]  = 1;
  ram[22573]  = 0;
  ram[22574]  = 0;
  ram[22575]  = 1;
  ram[22576]  = 1;
  ram[22577]  = 1;
  ram[22578]  = 1;
  ram[22579]  = 1;
  ram[22580]  = 0;
  ram[22581]  = 0;
  ram[22582]  = 0;
  ram[22583]  = 1;
  ram[22584]  = 1;
  ram[22585]  = 1;
  ram[22586]  = 1;
  ram[22587]  = 1;
  ram[22588]  = 1;
  ram[22589]  = 1;
  ram[22590]  = 1;
  ram[22591]  = 0;
  ram[22592]  = 1;
  ram[22593]  = 1;
  ram[22594]  = 1;
  ram[22595]  = 1;
  ram[22596]  = 1;
  ram[22597]  = 0;
  ram[22598]  = 1;
  ram[22599]  = 1;
  ram[22600]  = 1;
  ram[22601]  = 1;
  ram[22602]  = 1;
  ram[22603]  = 0;
  ram[22604]  = 1;
  ram[22605]  = 1;
  ram[22606]  = 0;
  ram[22607]  = 0;
  ram[22608]  = 1;
  ram[22609]  = 1;
  ram[22610]  = 1;
  ram[22611]  = 1;
  ram[22612]  = 1;
  ram[22613]  = 1;
  ram[22614]  = 1;
  ram[22615]  = 1;
  ram[22616]  = 1;
  ram[22617]  = 1;
  ram[22618]  = 1;
  ram[22619]  = 1;
  ram[22620]  = 1;
  ram[22621]  = 1;
  ram[22622]  = 0;
  ram[22623]  = 1;
  ram[22624]  = 1;
  ram[22625]  = 1;
  ram[22626]  = 1;
  ram[22627]  = 1;
  ram[22628]  = 0;
  ram[22629]  = 0;
  ram[22630]  = 1;
  ram[22631]  = 1;
  ram[22632]  = 0;
  ram[22633]  = 1;
  ram[22634]  = 1;
  ram[22635]  = 1;
  ram[22636]  = 1;
  ram[22637]  = 1;
  ram[22638]  = 0;
  ram[22639]  = 1;
  ram[22640]  = 1;
  ram[22641]  = 1;
  ram[22642]  = 0;
  ram[22643]  = 0;
  ram[22644]  = 1;
  ram[22645]  = 1;
  ram[22646]  = 1;
  ram[22647]  = 1;
  ram[22648]  = 0;
  ram[22649]  = 1;
  ram[22650]  = 1;
  ram[22651]  = 1;
  ram[22652]  = 1;
  ram[22653]  = 0;
  ram[22654]  = 0;
  ram[22655]  = 1;
  ram[22656]  = 1;
  ram[22657]  = 1;
  ram[22658]  = 1;
  ram[22659]  = 1;
  ram[22660]  = 1;
  ram[22661]  = 0;
  ram[22662]  = 1;
  ram[22663]  = 1;
  ram[22664]  = 0;
  ram[22665]  = 0;
  ram[22666]  = 1;
  ram[22667]  = 1;
  ram[22668]  = 1;
  ram[22669]  = 1;
  ram[22670]  = 1;
  ram[22671]  = 0;
  ram[22672]  = 1;
  ram[22673]  = 1;
  ram[22674]  = 1;
  ram[22675]  = 1;
  ram[22676]  = 1;
  ram[22677]  = 1;
  ram[22678]  = 1;
  ram[22679]  = 1;
  ram[22680]  = 0;
  ram[22681]  = 1;
  ram[22682]  = 1;
  ram[22683]  = 1;
  ram[22684]  = 1;
  ram[22685]  = 0;
  ram[22686]  = 1;
  ram[22687]  = 1;
  ram[22688]  = 1;
  ram[22689]  = 1;
  ram[22690]  = 1;
  ram[22691]  = 1;
  ram[22692]  = 1;
  ram[22693]  = 0;
  ram[22694]  = 1;
  ram[22695]  = 1;
  ram[22696]  = 1;
  ram[22697]  = 1;
  ram[22698]  = 1;
  ram[22699]  = 1;
  ram[22700]  = 1;
  ram[22701]  = 0;
  ram[22702]  = 0;
  ram[22703]  = 1;
  ram[22704]  = 1;
  ram[22705]  = 1;
  ram[22706]  = 1;
  ram[22707]  = 0;
  ram[22708]  = 1;
  ram[22709]  = 1;
  ram[22710]  = 1;
  ram[22711]  = 1;
  ram[22712]  = 1;
  ram[22713]  = 1;
  ram[22714]  = 1;
  ram[22715]  = 1;
  ram[22716]  = 1;
  ram[22717]  = 1;
  ram[22718]  = 1;
  ram[22719]  = 0;
  ram[22720]  = 0;
  ram[22721]  = 0;
  ram[22722]  = 1;
  ram[22723]  = 1;
  ram[22724]  = 1;
  ram[22725]  = 0;
  ram[22726]  = 1;
  ram[22727]  = 1;
  ram[22728]  = 1;
  ram[22729]  = 1;
  ram[22730]  = 1;
  ram[22731]  = 0;
  ram[22732]  = 1;
  ram[22733]  = 1;
  ram[22734]  = 1;
  ram[22735]  = 1;
  ram[22736]  = 0;
  ram[22737]  = 1;
  ram[22738]  = 1;
  ram[22739]  = 1;
  ram[22740]  = 0;
  ram[22741]  = 1;
  ram[22742]  = 1;
  ram[22743]  = 1;
  ram[22744]  = 1;
  ram[22745]  = 1;
  ram[22746]  = 0;
  ram[22747]  = 0;
  ram[22748]  = 1;
  ram[22749]  = 1;
  ram[22750]  = 1;
  ram[22751]  = 1;
  ram[22752]  = 1;
  ram[22753]  = 1;
  ram[22754]  = 1;
  ram[22755]  = 1;
  ram[22756]  = 1;
  ram[22757]  = 1;
  ram[22758]  = 1;
  ram[22759]  = 1;
  ram[22760]  = 1;
  ram[22761]  = 1;
  ram[22762]  = 1;
  ram[22763]  = 1;
  ram[22764]  = 1;
  ram[22765]  = 1;
  ram[22766]  = 1;
  ram[22767]  = 1;
  ram[22768]  = 1;
  ram[22769]  = 1;
  ram[22770]  = 1;
  ram[22771]  = 1;
  ram[22772]  = 1;
  ram[22773]  = 1;
  ram[22774]  = 1;
  ram[22775]  = 1;
  ram[22776]  = 1;
  ram[22777]  = 1;
  ram[22778]  = 1;
  ram[22779]  = 1;
  ram[22780]  = 1;
  ram[22781]  = 1;
  ram[22782]  = 1;
  ram[22783]  = 1;
  ram[22784]  = 1;
  ram[22785]  = 1;
  ram[22786]  = 1;
  ram[22787]  = 1;
  ram[22788]  = 1;
  ram[22789]  = 1;
  ram[22790]  = 1;
  ram[22791]  = 1;
  ram[22792]  = 1;
  ram[22793]  = 1;
  ram[22794]  = 1;
  ram[22795]  = 1;
  ram[22796]  = 1;
  ram[22797]  = 1;
  ram[22798]  = 1;
  ram[22799]  = 1;
  ram[22800]  = 1;
  ram[22801]  = 1;
  ram[22802]  = 1;
  ram[22803]  = 1;
  ram[22804]  = 1;
  ram[22805]  = 1;
  ram[22806]  = 1;
  ram[22807]  = 1;
  ram[22808]  = 1;
  ram[22809]  = 1;
  ram[22810]  = 1;
  ram[22811]  = 1;
  ram[22812]  = 1;
  ram[22813]  = 1;
  ram[22814]  = 1;
  ram[22815]  = 1;
  ram[22816]  = 1;
  ram[22817]  = 1;
  ram[22818]  = 1;
  ram[22819]  = 1;
  ram[22820]  = 1;
  ram[22821]  = 1;
  ram[22822]  = 1;
  ram[22823]  = 1;
  ram[22824]  = 1;
  ram[22825]  = 1;
  ram[22826]  = 1;
  ram[22827]  = 1;
  ram[22828]  = 1;
  ram[22829]  = 1;
  ram[22830]  = 1;
  ram[22831]  = 1;
  ram[22832]  = 1;
  ram[22833]  = 1;
  ram[22834]  = 1;
  ram[22835]  = 1;
  ram[22836]  = 1;
  ram[22837]  = 1;
  ram[22838]  = 1;
  ram[22839]  = 1;
  ram[22840]  = 1;
  ram[22841]  = 1;
  ram[22842]  = 1;
  ram[22843]  = 1;
  ram[22844]  = 1;
  ram[22845]  = 0;
  ram[22846]  = 1;
  ram[22847]  = 1;
  ram[22848]  = 1;
  ram[22849]  = 1;
  ram[22850]  = 1;
  ram[22851]  = 1;
  ram[22852]  = 1;
  ram[22853]  = 1;
  ram[22854]  = 1;
  ram[22855]  = 0;
  ram[22856]  = 1;
  ram[22857]  = 1;
  ram[22858]  = 1;
  ram[22859]  = 1;
  ram[22860]  = 1;
  ram[22861]  = 0;
  ram[22862]  = 1;
  ram[22863]  = 1;
  ram[22864]  = 1;
  ram[22865]  = 1;
  ram[22866]  = 1;
  ram[22867]  = 1;
  ram[22868]  = 1;
  ram[22869]  = 1;
  ram[22870]  = 1;
  ram[22871]  = 1;
  ram[22872]  = 1;
  ram[22873]  = 1;
  ram[22874]  = 0;
  ram[22875]  = 0;
  ram[22876]  = 1;
  ram[22877]  = 1;
  ram[22878]  = 1;
  ram[22879]  = 1;
  ram[22880]  = 1;
  ram[22881]  = 1;
  ram[22882]  = 0;
  ram[22883]  = 1;
  ram[22884]  = 1;
  ram[22885]  = 1;
  ram[22886]  = 1;
  ram[22887]  = 1;
  ram[22888]  = 1;
  ram[22889]  = 1;
  ram[22890]  = 1;
  ram[22891]  = 0;
  ram[22892]  = 1;
  ram[22893]  = 1;
  ram[22894]  = 1;
  ram[22895]  = 1;
  ram[22896]  = 1;
  ram[22897]  = 0;
  ram[22898]  = 1;
  ram[22899]  = 1;
  ram[22900]  = 1;
  ram[22901]  = 1;
  ram[22902]  = 1;
  ram[22903]  = 0;
  ram[22904]  = 1;
  ram[22905]  = 1;
  ram[22906]  = 0;
  ram[22907]  = 0;
  ram[22908]  = 1;
  ram[22909]  = 1;
  ram[22910]  = 1;
  ram[22911]  = 1;
  ram[22912]  = 1;
  ram[22913]  = 1;
  ram[22914]  = 1;
  ram[22915]  = 1;
  ram[22916]  = 1;
  ram[22917]  = 1;
  ram[22918]  = 1;
  ram[22919]  = 1;
  ram[22920]  = 1;
  ram[22921]  = 1;
  ram[22922]  = 0;
  ram[22923]  = 1;
  ram[22924]  = 1;
  ram[22925]  = 1;
  ram[22926]  = 1;
  ram[22927]  = 1;
  ram[22928]  = 1;
  ram[22929]  = 0;
  ram[22930]  = 1;
  ram[22931]  = 1;
  ram[22932]  = 0;
  ram[22933]  = 1;
  ram[22934]  = 1;
  ram[22935]  = 1;
  ram[22936]  = 1;
  ram[22937]  = 1;
  ram[22938]  = 0;
  ram[22939]  = 1;
  ram[22940]  = 1;
  ram[22941]  = 1;
  ram[22942]  = 0;
  ram[22943]  = 0;
  ram[22944]  = 1;
  ram[22945]  = 1;
  ram[22946]  = 1;
  ram[22947]  = 1;
  ram[22948]  = 0;
  ram[22949]  = 1;
  ram[22950]  = 1;
  ram[22951]  = 1;
  ram[22952]  = 1;
  ram[22953]  = 0;
  ram[22954]  = 0;
  ram[22955]  = 1;
  ram[22956]  = 1;
  ram[22957]  = 1;
  ram[22958]  = 1;
  ram[22959]  = 1;
  ram[22960]  = 1;
  ram[22961]  = 0;
  ram[22962]  = 1;
  ram[22963]  = 1;
  ram[22964]  = 0;
  ram[22965]  = 0;
  ram[22966]  = 1;
  ram[22967]  = 1;
  ram[22968]  = 1;
  ram[22969]  = 1;
  ram[22970]  = 1;
  ram[22971]  = 0;
  ram[22972]  = 1;
  ram[22973]  = 1;
  ram[22974]  = 1;
  ram[22975]  = 1;
  ram[22976]  = 1;
  ram[22977]  = 1;
  ram[22978]  = 1;
  ram[22979]  = 1;
  ram[22980]  = 0;
  ram[22981]  = 1;
  ram[22982]  = 1;
  ram[22983]  = 1;
  ram[22984]  = 1;
  ram[22985]  = 0;
  ram[22986]  = 1;
  ram[22987]  = 1;
  ram[22988]  = 1;
  ram[22989]  = 1;
  ram[22990]  = 1;
  ram[22991]  = 1;
  ram[22992]  = 1;
  ram[22993]  = 0;
  ram[22994]  = 1;
  ram[22995]  = 1;
  ram[22996]  = 1;
  ram[22997]  = 1;
  ram[22998]  = 1;
  ram[22999]  = 1;
  ram[23000]  = 1;
  ram[23001]  = 0;
  ram[23002]  = 0;
  ram[23003]  = 1;
  ram[23004]  = 1;
  ram[23005]  = 1;
  ram[23006]  = 1;
  ram[23007]  = 0;
  ram[23008]  = 1;
  ram[23009]  = 1;
  ram[23010]  = 1;
  ram[23011]  = 1;
  ram[23012]  = 1;
  ram[23013]  = 1;
  ram[23014]  = 1;
  ram[23015]  = 1;
  ram[23016]  = 1;
  ram[23017]  = 1;
  ram[23018]  = 1;
  ram[23019]  = 1;
  ram[23020]  = 1;
  ram[23021]  = 0;
  ram[23022]  = 1;
  ram[23023]  = 1;
  ram[23024]  = 1;
  ram[23025]  = 0;
  ram[23026]  = 1;
  ram[23027]  = 1;
  ram[23028]  = 1;
  ram[23029]  = 1;
  ram[23030]  = 0;
  ram[23031]  = 0;
  ram[23032]  = 1;
  ram[23033]  = 1;
  ram[23034]  = 1;
  ram[23035]  = 1;
  ram[23036]  = 0;
  ram[23037]  = 1;
  ram[23038]  = 1;
  ram[23039]  = 1;
  ram[23040]  = 0;
  ram[23041]  = 1;
  ram[23042]  = 1;
  ram[23043]  = 1;
  ram[23044]  = 1;
  ram[23045]  = 1;
  ram[23046]  = 0;
  ram[23047]  = 0;
  ram[23048]  = 1;
  ram[23049]  = 1;
  ram[23050]  = 1;
  ram[23051]  = 1;
  ram[23052]  = 1;
  ram[23053]  = 1;
  ram[23054]  = 1;
  ram[23055]  = 1;
  ram[23056]  = 1;
  ram[23057]  = 1;
  ram[23058]  = 1;
  ram[23059]  = 1;
  ram[23060]  = 1;
  ram[23061]  = 1;
  ram[23062]  = 1;
  ram[23063]  = 1;
  ram[23064]  = 1;
  ram[23065]  = 1;
  ram[23066]  = 1;
  ram[23067]  = 1;
  ram[23068]  = 1;
  ram[23069]  = 1;
  ram[23070]  = 1;
  ram[23071]  = 1;
  ram[23072]  = 1;
  ram[23073]  = 1;
  ram[23074]  = 1;
  ram[23075]  = 1;
  ram[23076]  = 1;
  ram[23077]  = 1;
  ram[23078]  = 1;
  ram[23079]  = 1;
  ram[23080]  = 1;
  ram[23081]  = 1;
  ram[23082]  = 1;
  ram[23083]  = 1;
  ram[23084]  = 1;
  ram[23085]  = 1;
  ram[23086]  = 1;
  ram[23087]  = 1;
  ram[23088]  = 1;
  ram[23089]  = 1;
  ram[23090]  = 1;
  ram[23091]  = 1;
  ram[23092]  = 1;
  ram[23093]  = 1;
  ram[23094]  = 1;
  ram[23095]  = 1;
  ram[23096]  = 1;
  ram[23097]  = 1;
  ram[23098]  = 1;
  ram[23099]  = 1;
  ram[23100]  = 1;
  ram[23101]  = 1;
  ram[23102]  = 1;
  ram[23103]  = 1;
  ram[23104]  = 1;
  ram[23105]  = 1;
  ram[23106]  = 1;
  ram[23107]  = 1;
  ram[23108]  = 1;
  ram[23109]  = 1;
  ram[23110]  = 1;
  ram[23111]  = 1;
  ram[23112]  = 1;
  ram[23113]  = 1;
  ram[23114]  = 1;
  ram[23115]  = 1;
  ram[23116]  = 1;
  ram[23117]  = 1;
  ram[23118]  = 1;
  ram[23119]  = 1;
  ram[23120]  = 1;
  ram[23121]  = 1;
  ram[23122]  = 1;
  ram[23123]  = 1;
  ram[23124]  = 1;
  ram[23125]  = 1;
  ram[23126]  = 1;
  ram[23127]  = 1;
  ram[23128]  = 1;
  ram[23129]  = 1;
  ram[23130]  = 1;
  ram[23131]  = 1;
  ram[23132]  = 1;
  ram[23133]  = 1;
  ram[23134]  = 1;
  ram[23135]  = 1;
  ram[23136]  = 1;
  ram[23137]  = 1;
  ram[23138]  = 1;
  ram[23139]  = 1;
  ram[23140]  = 1;
  ram[23141]  = 1;
  ram[23142]  = 1;
  ram[23143]  = 1;
  ram[23144]  = 1;
  ram[23145]  = 0;
  ram[23146]  = 1;
  ram[23147]  = 1;
  ram[23148]  = 1;
  ram[23149]  = 1;
  ram[23150]  = 1;
  ram[23151]  = 1;
  ram[23152]  = 1;
  ram[23153]  = 1;
  ram[23154]  = 1;
  ram[23155]  = 0;
  ram[23156]  = 1;
  ram[23157]  = 1;
  ram[23158]  = 1;
  ram[23159]  = 1;
  ram[23160]  = 1;
  ram[23161]  = 0;
  ram[23162]  = 1;
  ram[23163]  = 1;
  ram[23164]  = 1;
  ram[23165]  = 1;
  ram[23166]  = 1;
  ram[23167]  = 1;
  ram[23168]  = 1;
  ram[23169]  = 1;
  ram[23170]  = 1;
  ram[23171]  = 1;
  ram[23172]  = 1;
  ram[23173]  = 1;
  ram[23174]  = 1;
  ram[23175]  = 0;
  ram[23176]  = 1;
  ram[23177]  = 1;
  ram[23178]  = 1;
  ram[23179]  = 1;
  ram[23180]  = 1;
  ram[23181]  = 1;
  ram[23182]  = 0;
  ram[23183]  = 0;
  ram[23184]  = 1;
  ram[23185]  = 1;
  ram[23186]  = 1;
  ram[23187]  = 1;
  ram[23188]  = 1;
  ram[23189]  = 1;
  ram[23190]  = 1;
  ram[23191]  = 0;
  ram[23192]  = 1;
  ram[23193]  = 1;
  ram[23194]  = 1;
  ram[23195]  = 1;
  ram[23196]  = 1;
  ram[23197]  = 0;
  ram[23198]  = 1;
  ram[23199]  = 1;
  ram[23200]  = 1;
  ram[23201]  = 1;
  ram[23202]  = 1;
  ram[23203]  = 0;
  ram[23204]  = 1;
  ram[23205]  = 1;
  ram[23206]  = 0;
  ram[23207]  = 0;
  ram[23208]  = 1;
  ram[23209]  = 1;
  ram[23210]  = 1;
  ram[23211]  = 1;
  ram[23212]  = 1;
  ram[23213]  = 1;
  ram[23214]  = 1;
  ram[23215]  = 1;
  ram[23216]  = 1;
  ram[23217]  = 1;
  ram[23218]  = 1;
  ram[23219]  = 1;
  ram[23220]  = 1;
  ram[23221]  = 1;
  ram[23222]  = 0;
  ram[23223]  = 1;
  ram[23224]  = 1;
  ram[23225]  = 1;
  ram[23226]  = 1;
  ram[23227]  = 1;
  ram[23228]  = 0;
  ram[23229]  = 0;
  ram[23230]  = 1;
  ram[23231]  = 1;
  ram[23232]  = 0;
  ram[23233]  = 1;
  ram[23234]  = 1;
  ram[23235]  = 1;
  ram[23236]  = 1;
  ram[23237]  = 1;
  ram[23238]  = 0;
  ram[23239]  = 1;
  ram[23240]  = 1;
  ram[23241]  = 1;
  ram[23242]  = 0;
  ram[23243]  = 0;
  ram[23244]  = 1;
  ram[23245]  = 1;
  ram[23246]  = 1;
  ram[23247]  = 1;
  ram[23248]  = 0;
  ram[23249]  = 1;
  ram[23250]  = 1;
  ram[23251]  = 1;
  ram[23252]  = 1;
  ram[23253]  = 0;
  ram[23254]  = 0;
  ram[23255]  = 1;
  ram[23256]  = 1;
  ram[23257]  = 1;
  ram[23258]  = 1;
  ram[23259]  = 1;
  ram[23260]  = 1;
  ram[23261]  = 0;
  ram[23262]  = 1;
  ram[23263]  = 1;
  ram[23264]  = 0;
  ram[23265]  = 0;
  ram[23266]  = 1;
  ram[23267]  = 1;
  ram[23268]  = 1;
  ram[23269]  = 1;
  ram[23270]  = 1;
  ram[23271]  = 0;
  ram[23272]  = 1;
  ram[23273]  = 1;
  ram[23274]  = 1;
  ram[23275]  = 1;
  ram[23276]  = 1;
  ram[23277]  = 1;
  ram[23278]  = 1;
  ram[23279]  = 1;
  ram[23280]  = 0;
  ram[23281]  = 1;
  ram[23282]  = 1;
  ram[23283]  = 1;
  ram[23284]  = 1;
  ram[23285]  = 0;
  ram[23286]  = 1;
  ram[23287]  = 1;
  ram[23288]  = 1;
  ram[23289]  = 1;
  ram[23290]  = 1;
  ram[23291]  = 1;
  ram[23292]  = 1;
  ram[23293]  = 0;
  ram[23294]  = 1;
  ram[23295]  = 1;
  ram[23296]  = 1;
  ram[23297]  = 1;
  ram[23298]  = 1;
  ram[23299]  = 1;
  ram[23300]  = 1;
  ram[23301]  = 0;
  ram[23302]  = 0;
  ram[23303]  = 1;
  ram[23304]  = 1;
  ram[23305]  = 1;
  ram[23306]  = 1;
  ram[23307]  = 0;
  ram[23308]  = 1;
  ram[23309]  = 1;
  ram[23310]  = 1;
  ram[23311]  = 1;
  ram[23312]  = 1;
  ram[23313]  = 1;
  ram[23314]  = 1;
  ram[23315]  = 1;
  ram[23316]  = 1;
  ram[23317]  = 1;
  ram[23318]  = 1;
  ram[23319]  = 1;
  ram[23320]  = 1;
  ram[23321]  = 0;
  ram[23322]  = 0;
  ram[23323]  = 1;
  ram[23324]  = 1;
  ram[23325]  = 0;
  ram[23326]  = 1;
  ram[23327]  = 1;
  ram[23328]  = 1;
  ram[23329]  = 1;
  ram[23330]  = 0;
  ram[23331]  = 1;
  ram[23332]  = 1;
  ram[23333]  = 1;
  ram[23334]  = 1;
  ram[23335]  = 1;
  ram[23336]  = 0;
  ram[23337]  = 1;
  ram[23338]  = 1;
  ram[23339]  = 1;
  ram[23340]  = 0;
  ram[23341]  = 1;
  ram[23342]  = 1;
  ram[23343]  = 1;
  ram[23344]  = 1;
  ram[23345]  = 1;
  ram[23346]  = 0;
  ram[23347]  = 0;
  ram[23348]  = 1;
  ram[23349]  = 1;
  ram[23350]  = 1;
  ram[23351]  = 1;
  ram[23352]  = 1;
  ram[23353]  = 1;
  ram[23354]  = 1;
  ram[23355]  = 1;
  ram[23356]  = 1;
  ram[23357]  = 1;
  ram[23358]  = 1;
  ram[23359]  = 1;
  ram[23360]  = 1;
  ram[23361]  = 1;
  ram[23362]  = 1;
  ram[23363]  = 1;
  ram[23364]  = 1;
  ram[23365]  = 1;
  ram[23366]  = 1;
  ram[23367]  = 1;
  ram[23368]  = 1;
  ram[23369]  = 1;
  ram[23370]  = 1;
  ram[23371]  = 1;
  ram[23372]  = 1;
  ram[23373]  = 1;
  ram[23374]  = 1;
  ram[23375]  = 1;
  ram[23376]  = 1;
  ram[23377]  = 1;
  ram[23378]  = 1;
  ram[23379]  = 1;
  ram[23380]  = 1;
  ram[23381]  = 1;
  ram[23382]  = 1;
  ram[23383]  = 1;
  ram[23384]  = 1;
  ram[23385]  = 1;
  ram[23386]  = 1;
  ram[23387]  = 1;
  ram[23388]  = 1;
  ram[23389]  = 1;
  ram[23390]  = 1;
  ram[23391]  = 1;
  ram[23392]  = 1;
  ram[23393]  = 1;
  ram[23394]  = 1;
  ram[23395]  = 1;
  ram[23396]  = 1;
  ram[23397]  = 1;
  ram[23398]  = 1;
  ram[23399]  = 1;
  ram[23400]  = 1;
  ram[23401]  = 1;
  ram[23402]  = 1;
  ram[23403]  = 1;
  ram[23404]  = 1;
  ram[23405]  = 1;
  ram[23406]  = 1;
  ram[23407]  = 1;
  ram[23408]  = 1;
  ram[23409]  = 1;
  ram[23410]  = 1;
  ram[23411]  = 1;
  ram[23412]  = 1;
  ram[23413]  = 1;
  ram[23414]  = 1;
  ram[23415]  = 1;
  ram[23416]  = 1;
  ram[23417]  = 1;
  ram[23418]  = 1;
  ram[23419]  = 1;
  ram[23420]  = 1;
  ram[23421]  = 1;
  ram[23422]  = 1;
  ram[23423]  = 1;
  ram[23424]  = 1;
  ram[23425]  = 1;
  ram[23426]  = 1;
  ram[23427]  = 1;
  ram[23428]  = 1;
  ram[23429]  = 1;
  ram[23430]  = 1;
  ram[23431]  = 1;
  ram[23432]  = 1;
  ram[23433]  = 1;
  ram[23434]  = 1;
  ram[23435]  = 1;
  ram[23436]  = 1;
  ram[23437]  = 1;
  ram[23438]  = 1;
  ram[23439]  = 1;
  ram[23440]  = 1;
  ram[23441]  = 1;
  ram[23442]  = 1;
  ram[23443]  = 1;
  ram[23444]  = 1;
  ram[23445]  = 0;
  ram[23446]  = 1;
  ram[23447]  = 1;
  ram[23448]  = 1;
  ram[23449]  = 1;
  ram[23450]  = 1;
  ram[23451]  = 1;
  ram[23452]  = 1;
  ram[23453]  = 1;
  ram[23454]  = 1;
  ram[23455]  = 0;
  ram[23456]  = 1;
  ram[23457]  = 1;
  ram[23458]  = 1;
  ram[23459]  = 1;
  ram[23460]  = 1;
  ram[23461]  = 0;
  ram[23462]  = 1;
  ram[23463]  = 1;
  ram[23464]  = 1;
  ram[23465]  = 1;
  ram[23466]  = 1;
  ram[23467]  = 1;
  ram[23468]  = 1;
  ram[23469]  = 1;
  ram[23470]  = 1;
  ram[23471]  = 1;
  ram[23472]  = 1;
  ram[23473]  = 1;
  ram[23474]  = 1;
  ram[23475]  = 0;
  ram[23476]  = 1;
  ram[23477]  = 1;
  ram[23478]  = 1;
  ram[23479]  = 1;
  ram[23480]  = 1;
  ram[23481]  = 1;
  ram[23482]  = 0;
  ram[23483]  = 0;
  ram[23484]  = 1;
  ram[23485]  = 1;
  ram[23486]  = 1;
  ram[23487]  = 1;
  ram[23488]  = 1;
  ram[23489]  = 1;
  ram[23490]  = 1;
  ram[23491]  = 0;
  ram[23492]  = 1;
  ram[23493]  = 1;
  ram[23494]  = 1;
  ram[23495]  = 1;
  ram[23496]  = 1;
  ram[23497]  = 0;
  ram[23498]  = 1;
  ram[23499]  = 1;
  ram[23500]  = 1;
  ram[23501]  = 1;
  ram[23502]  = 1;
  ram[23503]  = 0;
  ram[23504]  = 1;
  ram[23505]  = 1;
  ram[23506]  = 1;
  ram[23507]  = 0;
  ram[23508]  = 1;
  ram[23509]  = 1;
  ram[23510]  = 1;
  ram[23511]  = 1;
  ram[23512]  = 1;
  ram[23513]  = 1;
  ram[23514]  = 1;
  ram[23515]  = 1;
  ram[23516]  = 1;
  ram[23517]  = 1;
  ram[23518]  = 1;
  ram[23519]  = 1;
  ram[23520]  = 1;
  ram[23521]  = 1;
  ram[23522]  = 0;
  ram[23523]  = 1;
  ram[23524]  = 1;
  ram[23525]  = 1;
  ram[23526]  = 1;
  ram[23527]  = 1;
  ram[23528]  = 0;
  ram[23529]  = 0;
  ram[23530]  = 1;
  ram[23531]  = 1;
  ram[23532]  = 0;
  ram[23533]  = 1;
  ram[23534]  = 1;
  ram[23535]  = 1;
  ram[23536]  = 1;
  ram[23537]  = 1;
  ram[23538]  = 0;
  ram[23539]  = 1;
  ram[23540]  = 1;
  ram[23541]  = 1;
  ram[23542]  = 0;
  ram[23543]  = 0;
  ram[23544]  = 1;
  ram[23545]  = 1;
  ram[23546]  = 1;
  ram[23547]  = 1;
  ram[23548]  = 0;
  ram[23549]  = 1;
  ram[23550]  = 1;
  ram[23551]  = 1;
  ram[23552]  = 1;
  ram[23553]  = 1;
  ram[23554]  = 0;
  ram[23555]  = 1;
  ram[23556]  = 1;
  ram[23557]  = 1;
  ram[23558]  = 1;
  ram[23559]  = 1;
  ram[23560]  = 1;
  ram[23561]  = 0;
  ram[23562]  = 1;
  ram[23563]  = 1;
  ram[23564]  = 0;
  ram[23565]  = 0;
  ram[23566]  = 1;
  ram[23567]  = 1;
  ram[23568]  = 1;
  ram[23569]  = 1;
  ram[23570]  = 1;
  ram[23571]  = 0;
  ram[23572]  = 1;
  ram[23573]  = 1;
  ram[23574]  = 1;
  ram[23575]  = 1;
  ram[23576]  = 1;
  ram[23577]  = 1;
  ram[23578]  = 1;
  ram[23579]  = 1;
  ram[23580]  = 0;
  ram[23581]  = 1;
  ram[23582]  = 1;
  ram[23583]  = 1;
  ram[23584]  = 1;
  ram[23585]  = 0;
  ram[23586]  = 0;
  ram[23587]  = 1;
  ram[23588]  = 1;
  ram[23589]  = 1;
  ram[23590]  = 1;
  ram[23591]  = 1;
  ram[23592]  = 0;
  ram[23593]  = 0;
  ram[23594]  = 1;
  ram[23595]  = 1;
  ram[23596]  = 1;
  ram[23597]  = 1;
  ram[23598]  = 1;
  ram[23599]  = 1;
  ram[23600]  = 1;
  ram[23601]  = 0;
  ram[23602]  = 0;
  ram[23603]  = 1;
  ram[23604]  = 1;
  ram[23605]  = 1;
  ram[23606]  = 1;
  ram[23607]  = 0;
  ram[23608]  = 0;
  ram[23609]  = 1;
  ram[23610]  = 1;
  ram[23611]  = 1;
  ram[23612]  = 1;
  ram[23613]  = 1;
  ram[23614]  = 1;
  ram[23615]  = 1;
  ram[23616]  = 1;
  ram[23617]  = 1;
  ram[23618]  = 1;
  ram[23619]  = 1;
  ram[23620]  = 1;
  ram[23621]  = 1;
  ram[23622]  = 0;
  ram[23623]  = 1;
  ram[23624]  = 1;
  ram[23625]  = 0;
  ram[23626]  = 1;
  ram[23627]  = 1;
  ram[23628]  = 1;
  ram[23629]  = 1;
  ram[23630]  = 0;
  ram[23631]  = 1;
  ram[23632]  = 1;
  ram[23633]  = 1;
  ram[23634]  = 1;
  ram[23635]  = 1;
  ram[23636]  = 0;
  ram[23637]  = 1;
  ram[23638]  = 1;
  ram[23639]  = 1;
  ram[23640]  = 0;
  ram[23641]  = 1;
  ram[23642]  = 1;
  ram[23643]  = 1;
  ram[23644]  = 1;
  ram[23645]  = 1;
  ram[23646]  = 0;
  ram[23647]  = 0;
  ram[23648]  = 1;
  ram[23649]  = 1;
  ram[23650]  = 1;
  ram[23651]  = 1;
  ram[23652]  = 1;
  ram[23653]  = 1;
  ram[23654]  = 1;
  ram[23655]  = 1;
  ram[23656]  = 1;
  ram[23657]  = 1;
  ram[23658]  = 1;
  ram[23659]  = 1;
  ram[23660]  = 1;
  ram[23661]  = 1;
  ram[23662]  = 1;
  ram[23663]  = 1;
  ram[23664]  = 1;
  ram[23665]  = 1;
  ram[23666]  = 1;
  ram[23667]  = 1;
  ram[23668]  = 1;
  ram[23669]  = 1;
  ram[23670]  = 1;
  ram[23671]  = 1;
  ram[23672]  = 1;
  ram[23673]  = 1;
  ram[23674]  = 1;
  ram[23675]  = 1;
  ram[23676]  = 1;
  ram[23677]  = 1;
  ram[23678]  = 1;
  ram[23679]  = 1;
  ram[23680]  = 1;
  ram[23681]  = 1;
  ram[23682]  = 1;
  ram[23683]  = 1;
  ram[23684]  = 1;
  ram[23685]  = 1;
  ram[23686]  = 1;
  ram[23687]  = 1;
  ram[23688]  = 1;
  ram[23689]  = 1;
  ram[23690]  = 1;
  ram[23691]  = 1;
  ram[23692]  = 1;
  ram[23693]  = 1;
  ram[23694]  = 1;
  ram[23695]  = 1;
  ram[23696]  = 1;
  ram[23697]  = 1;
  ram[23698]  = 1;
  ram[23699]  = 1;
  ram[23700]  = 1;
  ram[23701]  = 1;
  ram[23702]  = 1;
  ram[23703]  = 1;
  ram[23704]  = 1;
  ram[23705]  = 1;
  ram[23706]  = 1;
  ram[23707]  = 1;
  ram[23708]  = 1;
  ram[23709]  = 1;
  ram[23710]  = 1;
  ram[23711]  = 1;
  ram[23712]  = 1;
  ram[23713]  = 1;
  ram[23714]  = 1;
  ram[23715]  = 1;
  ram[23716]  = 1;
  ram[23717]  = 1;
  ram[23718]  = 1;
  ram[23719]  = 1;
  ram[23720]  = 1;
  ram[23721]  = 1;
  ram[23722]  = 1;
  ram[23723]  = 1;
  ram[23724]  = 1;
  ram[23725]  = 1;
  ram[23726]  = 1;
  ram[23727]  = 1;
  ram[23728]  = 1;
  ram[23729]  = 1;
  ram[23730]  = 1;
  ram[23731]  = 1;
  ram[23732]  = 1;
  ram[23733]  = 1;
  ram[23734]  = 1;
  ram[23735]  = 1;
  ram[23736]  = 1;
  ram[23737]  = 1;
  ram[23738]  = 1;
  ram[23739]  = 1;
  ram[23740]  = 1;
  ram[23741]  = 1;
  ram[23742]  = 1;
  ram[23743]  = 1;
  ram[23744]  = 1;
  ram[23745]  = 0;
  ram[23746]  = 1;
  ram[23747]  = 1;
  ram[23748]  = 1;
  ram[23749]  = 1;
  ram[23750]  = 1;
  ram[23751]  = 1;
  ram[23752]  = 1;
  ram[23753]  = 1;
  ram[23754]  = 1;
  ram[23755]  = 0;
  ram[23756]  = 1;
  ram[23757]  = 1;
  ram[23758]  = 1;
  ram[23759]  = 1;
  ram[23760]  = 1;
  ram[23761]  = 0;
  ram[23762]  = 1;
  ram[23763]  = 1;
  ram[23764]  = 1;
  ram[23765]  = 1;
  ram[23766]  = 1;
  ram[23767]  = 0;
  ram[23768]  = 1;
  ram[23769]  = 1;
  ram[23770]  = 0;
  ram[23771]  = 1;
  ram[23772]  = 1;
  ram[23773]  = 1;
  ram[23774]  = 1;
  ram[23775]  = 0;
  ram[23776]  = 1;
  ram[23777]  = 0;
  ram[23778]  = 1;
  ram[23779]  = 1;
  ram[23780]  = 1;
  ram[23781]  = 1;
  ram[23782]  = 0;
  ram[23783]  = 0;
  ram[23784]  = 1;
  ram[23785]  = 1;
  ram[23786]  = 1;
  ram[23787]  = 1;
  ram[23788]  = 1;
  ram[23789]  = 1;
  ram[23790]  = 1;
  ram[23791]  = 0;
  ram[23792]  = 1;
  ram[23793]  = 1;
  ram[23794]  = 1;
  ram[23795]  = 1;
  ram[23796]  = 1;
  ram[23797]  = 0;
  ram[23798]  = 1;
  ram[23799]  = 1;
  ram[23800]  = 1;
  ram[23801]  = 1;
  ram[23802]  = 1;
  ram[23803]  = 0;
  ram[23804]  = 1;
  ram[23805]  = 1;
  ram[23806]  = 1;
  ram[23807]  = 0;
  ram[23808]  = 1;
  ram[23809]  = 1;
  ram[23810]  = 1;
  ram[23811]  = 1;
  ram[23812]  = 1;
  ram[23813]  = 0;
  ram[23814]  = 1;
  ram[23815]  = 1;
  ram[23816]  = 1;
  ram[23817]  = 1;
  ram[23818]  = 1;
  ram[23819]  = 1;
  ram[23820]  = 1;
  ram[23821]  = 1;
  ram[23822]  = 0;
  ram[23823]  = 1;
  ram[23824]  = 1;
  ram[23825]  = 1;
  ram[23826]  = 1;
  ram[23827]  = 1;
  ram[23828]  = 0;
  ram[23829]  = 1;
  ram[23830]  = 1;
  ram[23831]  = 1;
  ram[23832]  = 0;
  ram[23833]  = 1;
  ram[23834]  = 1;
  ram[23835]  = 1;
  ram[23836]  = 1;
  ram[23837]  = 0;
  ram[23838]  = 0;
  ram[23839]  = 1;
  ram[23840]  = 1;
  ram[23841]  = 1;
  ram[23842]  = 0;
  ram[23843]  = 0;
  ram[23844]  = 1;
  ram[23845]  = 1;
  ram[23846]  = 1;
  ram[23847]  = 1;
  ram[23848]  = 0;
  ram[23849]  = 1;
  ram[23850]  = 1;
  ram[23851]  = 1;
  ram[23852]  = 1;
  ram[23853]  = 1;
  ram[23854]  = 0;
  ram[23855]  = 1;
  ram[23856]  = 1;
  ram[23857]  = 1;
  ram[23858]  = 1;
  ram[23859]  = 1;
  ram[23860]  = 0;
  ram[23861]  = 0;
  ram[23862]  = 1;
  ram[23863]  = 1;
  ram[23864]  = 0;
  ram[23865]  = 0;
  ram[23866]  = 1;
  ram[23867]  = 1;
  ram[23868]  = 1;
  ram[23869]  = 1;
  ram[23870]  = 1;
  ram[23871]  = 0;
  ram[23872]  = 1;
  ram[23873]  = 1;
  ram[23874]  = 1;
  ram[23875]  = 1;
  ram[23876]  = 1;
  ram[23877]  = 1;
  ram[23878]  = 1;
  ram[23879]  = 1;
  ram[23880]  = 0;
  ram[23881]  = 1;
  ram[23882]  = 1;
  ram[23883]  = 1;
  ram[23884]  = 1;
  ram[23885]  = 1;
  ram[23886]  = 0;
  ram[23887]  = 1;
  ram[23888]  = 1;
  ram[23889]  = 1;
  ram[23890]  = 1;
  ram[23891]  = 1;
  ram[23892]  = 0;
  ram[23893]  = 1;
  ram[23894]  = 1;
  ram[23895]  = 1;
  ram[23896]  = 1;
  ram[23897]  = 1;
  ram[23898]  = 1;
  ram[23899]  = 1;
  ram[23900]  = 1;
  ram[23901]  = 0;
  ram[23902]  = 0;
  ram[23903]  = 1;
  ram[23904]  = 1;
  ram[23905]  = 1;
  ram[23906]  = 1;
  ram[23907]  = 0;
  ram[23908]  = 0;
  ram[23909]  = 1;
  ram[23910]  = 1;
  ram[23911]  = 1;
  ram[23912]  = 1;
  ram[23913]  = 1;
  ram[23914]  = 0;
  ram[23915]  = 1;
  ram[23916]  = 0;
  ram[23917]  = 1;
  ram[23918]  = 1;
  ram[23919]  = 1;
  ram[23920]  = 1;
  ram[23921]  = 1;
  ram[23922]  = 0;
  ram[23923]  = 1;
  ram[23924]  = 1;
  ram[23925]  = 0;
  ram[23926]  = 1;
  ram[23927]  = 1;
  ram[23928]  = 1;
  ram[23929]  = 1;
  ram[23930]  = 0;
  ram[23931]  = 1;
  ram[23932]  = 1;
  ram[23933]  = 1;
  ram[23934]  = 1;
  ram[23935]  = 0;
  ram[23936]  = 0;
  ram[23937]  = 1;
  ram[23938]  = 1;
  ram[23939]  = 1;
  ram[23940]  = 0;
  ram[23941]  = 1;
  ram[23942]  = 1;
  ram[23943]  = 1;
  ram[23944]  = 1;
  ram[23945]  = 1;
  ram[23946]  = 0;
  ram[23947]  = 0;
  ram[23948]  = 1;
  ram[23949]  = 1;
  ram[23950]  = 1;
  ram[23951]  = 1;
  ram[23952]  = 1;
  ram[23953]  = 1;
  ram[23954]  = 1;
  ram[23955]  = 1;
  ram[23956]  = 1;
  ram[23957]  = 1;
  ram[23958]  = 1;
  ram[23959]  = 1;
  ram[23960]  = 1;
  ram[23961]  = 1;
  ram[23962]  = 1;
  ram[23963]  = 1;
  ram[23964]  = 1;
  ram[23965]  = 1;
  ram[23966]  = 1;
  ram[23967]  = 1;
  ram[23968]  = 1;
  ram[23969]  = 1;
  ram[23970]  = 1;
  ram[23971]  = 1;
  ram[23972]  = 1;
  ram[23973]  = 1;
  ram[23974]  = 1;
  ram[23975]  = 1;
  ram[23976]  = 1;
  ram[23977]  = 1;
  ram[23978]  = 1;
  ram[23979]  = 1;
  ram[23980]  = 1;
  ram[23981]  = 1;
  ram[23982]  = 1;
  ram[23983]  = 1;
  ram[23984]  = 1;
  ram[23985]  = 1;
  ram[23986]  = 1;
  ram[23987]  = 1;
  ram[23988]  = 1;
  ram[23989]  = 1;
  ram[23990]  = 1;
  ram[23991]  = 1;
  ram[23992]  = 1;
  ram[23993]  = 1;
  ram[23994]  = 1;
  ram[23995]  = 1;
  ram[23996]  = 1;
  ram[23997]  = 1;
  ram[23998]  = 1;
  ram[23999]  = 1;
  ram[24000]  = 1;
  ram[24001]  = 1;
  ram[24002]  = 1;
  ram[24003]  = 1;
  ram[24004]  = 1;
  ram[24005]  = 1;
  ram[24006]  = 1;
  ram[24007]  = 1;
  ram[24008]  = 1;
  ram[24009]  = 1;
  ram[24010]  = 1;
  ram[24011]  = 1;
  ram[24012]  = 1;
  ram[24013]  = 1;
  ram[24014]  = 1;
  ram[24015]  = 1;
  ram[24016]  = 1;
  ram[24017]  = 1;
  ram[24018]  = 1;
  ram[24019]  = 1;
  ram[24020]  = 1;
  ram[24021]  = 1;
  ram[24022]  = 1;
  ram[24023]  = 1;
  ram[24024]  = 1;
  ram[24025]  = 1;
  ram[24026]  = 1;
  ram[24027]  = 1;
  ram[24028]  = 1;
  ram[24029]  = 1;
  ram[24030]  = 1;
  ram[24031]  = 1;
  ram[24032]  = 1;
  ram[24033]  = 1;
  ram[24034]  = 1;
  ram[24035]  = 1;
  ram[24036]  = 1;
  ram[24037]  = 1;
  ram[24038]  = 1;
  ram[24039]  = 1;
  ram[24040]  = 1;
  ram[24041]  = 1;
  ram[24042]  = 1;
  ram[24043]  = 1;
  ram[24044]  = 1;
  ram[24045]  = 0;
  ram[24046]  = 1;
  ram[24047]  = 1;
  ram[24048]  = 1;
  ram[24049]  = 1;
  ram[24050]  = 1;
  ram[24051]  = 1;
  ram[24052]  = 1;
  ram[24053]  = 1;
  ram[24054]  = 1;
  ram[24055]  = 0;
  ram[24056]  = 1;
  ram[24057]  = 1;
  ram[24058]  = 1;
  ram[24059]  = 1;
  ram[24060]  = 1;
  ram[24061]  = 0;
  ram[24062]  = 0;
  ram[24063]  = 1;
  ram[24064]  = 1;
  ram[24065]  = 1;
  ram[24066]  = 1;
  ram[24067]  = 0;
  ram[24068]  = 1;
  ram[24069]  = 1;
  ram[24070]  = 0;
  ram[24071]  = 1;
  ram[24072]  = 1;
  ram[24073]  = 1;
  ram[24074]  = 1;
  ram[24075]  = 0;
  ram[24076]  = 1;
  ram[24077]  = 0;
  ram[24078]  = 1;
  ram[24079]  = 1;
  ram[24080]  = 1;
  ram[24081]  = 1;
  ram[24082]  = 0;
  ram[24083]  = 0;
  ram[24084]  = 1;
  ram[24085]  = 1;
  ram[24086]  = 1;
  ram[24087]  = 1;
  ram[24088]  = 1;
  ram[24089]  = 1;
  ram[24090]  = 1;
  ram[24091]  = 0;
  ram[24092]  = 1;
  ram[24093]  = 1;
  ram[24094]  = 1;
  ram[24095]  = 1;
  ram[24096]  = 1;
  ram[24097]  = 0;
  ram[24098]  = 1;
  ram[24099]  = 1;
  ram[24100]  = 1;
  ram[24101]  = 1;
  ram[24102]  = 1;
  ram[24103]  = 0;
  ram[24104]  = 1;
  ram[24105]  = 1;
  ram[24106]  = 1;
  ram[24107]  = 0;
  ram[24108]  = 0;
  ram[24109]  = 1;
  ram[24110]  = 1;
  ram[24111]  = 1;
  ram[24112]  = 0;
  ram[24113]  = 0;
  ram[24114]  = 1;
  ram[24115]  = 1;
  ram[24116]  = 1;
  ram[24117]  = 1;
  ram[24118]  = 1;
  ram[24119]  = 1;
  ram[24120]  = 1;
  ram[24121]  = 1;
  ram[24122]  = 0;
  ram[24123]  = 1;
  ram[24124]  = 1;
  ram[24125]  = 1;
  ram[24126]  = 1;
  ram[24127]  = 0;
  ram[24128]  = 0;
  ram[24129]  = 1;
  ram[24130]  = 1;
  ram[24131]  = 1;
  ram[24132]  = 0;
  ram[24133]  = 1;
  ram[24134]  = 1;
  ram[24135]  = 1;
  ram[24136]  = 1;
  ram[24137]  = 0;
  ram[24138]  = 0;
  ram[24139]  = 1;
  ram[24140]  = 1;
  ram[24141]  = 1;
  ram[24142]  = 0;
  ram[24143]  = 0;
  ram[24144]  = 1;
  ram[24145]  = 1;
  ram[24146]  = 1;
  ram[24147]  = 1;
  ram[24148]  = 0;
  ram[24149]  = 1;
  ram[24150]  = 1;
  ram[24151]  = 1;
  ram[24152]  = 1;
  ram[24153]  = 1;
  ram[24154]  = 0;
  ram[24155]  = 0;
  ram[24156]  = 1;
  ram[24157]  = 1;
  ram[24158]  = 1;
  ram[24159]  = 1;
  ram[24160]  = 0;
  ram[24161]  = 1;
  ram[24162]  = 1;
  ram[24163]  = 1;
  ram[24164]  = 0;
  ram[24165]  = 0;
  ram[24166]  = 1;
  ram[24167]  = 1;
  ram[24168]  = 1;
  ram[24169]  = 1;
  ram[24170]  = 1;
  ram[24171]  = 0;
  ram[24172]  = 1;
  ram[24173]  = 1;
  ram[24174]  = 1;
  ram[24175]  = 1;
  ram[24176]  = 1;
  ram[24177]  = 1;
  ram[24178]  = 1;
  ram[24179]  = 1;
  ram[24180]  = 0;
  ram[24181]  = 1;
  ram[24182]  = 1;
  ram[24183]  = 1;
  ram[24184]  = 1;
  ram[24185]  = 1;
  ram[24186]  = 0;
  ram[24187]  = 1;
  ram[24188]  = 1;
  ram[24189]  = 1;
  ram[24190]  = 1;
  ram[24191]  = 1;
  ram[24192]  = 0;
  ram[24193]  = 1;
  ram[24194]  = 1;
  ram[24195]  = 1;
  ram[24196]  = 1;
  ram[24197]  = 1;
  ram[24198]  = 1;
  ram[24199]  = 1;
  ram[24200]  = 1;
  ram[24201]  = 0;
  ram[24202]  = 0;
  ram[24203]  = 1;
  ram[24204]  = 1;
  ram[24205]  = 1;
  ram[24206]  = 1;
  ram[24207]  = 1;
  ram[24208]  = 0;
  ram[24209]  = 1;
  ram[24210]  = 1;
  ram[24211]  = 1;
  ram[24212]  = 1;
  ram[24213]  = 0;
  ram[24214]  = 1;
  ram[24215]  = 1;
  ram[24216]  = 0;
  ram[24217]  = 1;
  ram[24218]  = 1;
  ram[24219]  = 1;
  ram[24220]  = 1;
  ram[24221]  = 0;
  ram[24222]  = 0;
  ram[24223]  = 1;
  ram[24224]  = 1;
  ram[24225]  = 0;
  ram[24226]  = 1;
  ram[24227]  = 1;
  ram[24228]  = 1;
  ram[24229]  = 1;
  ram[24230]  = 0;
  ram[24231]  = 1;
  ram[24232]  = 1;
  ram[24233]  = 1;
  ram[24234]  = 1;
  ram[24235]  = 0;
  ram[24236]  = 0;
  ram[24237]  = 1;
  ram[24238]  = 1;
  ram[24239]  = 1;
  ram[24240]  = 0;
  ram[24241]  = 1;
  ram[24242]  = 1;
  ram[24243]  = 1;
  ram[24244]  = 1;
  ram[24245]  = 1;
  ram[24246]  = 0;
  ram[24247]  = 0;
  ram[24248]  = 1;
  ram[24249]  = 1;
  ram[24250]  = 1;
  ram[24251]  = 1;
  ram[24252]  = 1;
  ram[24253]  = 1;
  ram[24254]  = 1;
  ram[24255]  = 1;
  ram[24256]  = 1;
  ram[24257]  = 1;
  ram[24258]  = 1;
  ram[24259]  = 1;
  ram[24260]  = 1;
  ram[24261]  = 1;
  ram[24262]  = 1;
  ram[24263]  = 1;
  ram[24264]  = 1;
  ram[24265]  = 1;
  ram[24266]  = 1;
  ram[24267]  = 1;
  ram[24268]  = 1;
  ram[24269]  = 1;
  ram[24270]  = 1;
  ram[24271]  = 1;
  ram[24272]  = 1;
  ram[24273]  = 1;
  ram[24274]  = 1;
  ram[24275]  = 1;
  ram[24276]  = 1;
  ram[24277]  = 1;
  ram[24278]  = 1;
  ram[24279]  = 1;
  ram[24280]  = 1;
  ram[24281]  = 1;
  ram[24282]  = 1;
  ram[24283]  = 1;
  ram[24284]  = 1;
  ram[24285]  = 1;
  ram[24286]  = 1;
  ram[24287]  = 1;
  ram[24288]  = 1;
  ram[24289]  = 1;
  ram[24290]  = 1;
  ram[24291]  = 1;
  ram[24292]  = 1;
  ram[24293]  = 1;
  ram[24294]  = 1;
  ram[24295]  = 1;
  ram[24296]  = 1;
  ram[24297]  = 1;
  ram[24298]  = 1;
  ram[24299]  = 1;
  ram[24300]  = 1;
  ram[24301]  = 1;
  ram[24302]  = 1;
  ram[24303]  = 1;
  ram[24304]  = 1;
  ram[24305]  = 1;
  ram[24306]  = 1;
  ram[24307]  = 1;
  ram[24308]  = 1;
  ram[24309]  = 1;
  ram[24310]  = 1;
  ram[24311]  = 1;
  ram[24312]  = 1;
  ram[24313]  = 1;
  ram[24314]  = 1;
  ram[24315]  = 1;
  ram[24316]  = 1;
  ram[24317]  = 1;
  ram[24318]  = 1;
  ram[24319]  = 1;
  ram[24320]  = 1;
  ram[24321]  = 1;
  ram[24322]  = 1;
  ram[24323]  = 1;
  ram[24324]  = 1;
  ram[24325]  = 1;
  ram[24326]  = 1;
  ram[24327]  = 1;
  ram[24328]  = 1;
  ram[24329]  = 1;
  ram[24330]  = 1;
  ram[24331]  = 1;
  ram[24332]  = 1;
  ram[24333]  = 1;
  ram[24334]  = 1;
  ram[24335]  = 1;
  ram[24336]  = 1;
  ram[24337]  = 1;
  ram[24338]  = 1;
  ram[24339]  = 1;
  ram[24340]  = 1;
  ram[24341]  = 1;
  ram[24342]  = 1;
  ram[24343]  = 1;
  ram[24344]  = 1;
  ram[24345]  = 0;
  ram[24346]  = 1;
  ram[24347]  = 1;
  ram[24348]  = 1;
  ram[24349]  = 1;
  ram[24350]  = 1;
  ram[24351]  = 1;
  ram[24352]  = 1;
  ram[24353]  = 1;
  ram[24354]  = 1;
  ram[24355]  = 0;
  ram[24356]  = 1;
  ram[24357]  = 1;
  ram[24358]  = 1;
  ram[24359]  = 1;
  ram[24360]  = 1;
  ram[24361]  = 1;
  ram[24362]  = 0;
  ram[24363]  = 0;
  ram[24364]  = 1;
  ram[24365]  = 1;
  ram[24366]  = 0;
  ram[24367]  = 0;
  ram[24368]  = 1;
  ram[24369]  = 1;
  ram[24370]  = 0;
  ram[24371]  = 0;
  ram[24372]  = 1;
  ram[24373]  = 1;
  ram[24374]  = 0;
  ram[24375]  = 0;
  ram[24376]  = 1;
  ram[24377]  = 1;
  ram[24378]  = 0;
  ram[24379]  = 1;
  ram[24380]  = 1;
  ram[24381]  = 1;
  ram[24382]  = 0;
  ram[24383]  = 1;
  ram[24384]  = 1;
  ram[24385]  = 1;
  ram[24386]  = 1;
  ram[24387]  = 1;
  ram[24388]  = 1;
  ram[24389]  = 1;
  ram[24390]  = 1;
  ram[24391]  = 0;
  ram[24392]  = 0;
  ram[24393]  = 1;
  ram[24394]  = 1;
  ram[24395]  = 1;
  ram[24396]  = 1;
  ram[24397]  = 0;
  ram[24398]  = 1;
  ram[24399]  = 1;
  ram[24400]  = 1;
  ram[24401]  = 1;
  ram[24402]  = 1;
  ram[24403]  = 0;
  ram[24404]  = 1;
  ram[24405]  = 1;
  ram[24406]  = 1;
  ram[24407]  = 1;
  ram[24408]  = 0;
  ram[24409]  = 0;
  ram[24410]  = 1;
  ram[24411]  = 0;
  ram[24412]  = 0;
  ram[24413]  = 1;
  ram[24414]  = 1;
  ram[24415]  = 1;
  ram[24416]  = 1;
  ram[24417]  = 1;
  ram[24418]  = 1;
  ram[24419]  = 1;
  ram[24420]  = 1;
  ram[24421]  = 1;
  ram[24422]  = 0;
  ram[24423]  = 0;
  ram[24424]  = 0;
  ram[24425]  = 0;
  ram[24426]  = 0;
  ram[24427]  = 0;
  ram[24428]  = 0;
  ram[24429]  = 1;
  ram[24430]  = 1;
  ram[24431]  = 1;
  ram[24432]  = 0;
  ram[24433]  = 0;
  ram[24434]  = 1;
  ram[24435]  = 1;
  ram[24436]  = 0;
  ram[24437]  = 1;
  ram[24438]  = 0;
  ram[24439]  = 1;
  ram[24440]  = 1;
  ram[24441]  = 1;
  ram[24442]  = 1;
  ram[24443]  = 0;
  ram[24444]  = 1;
  ram[24445]  = 1;
  ram[24446]  = 1;
  ram[24447]  = 1;
  ram[24448]  = 0;
  ram[24449]  = 0;
  ram[24450]  = 1;
  ram[24451]  = 1;
  ram[24452]  = 1;
  ram[24453]  = 1;
  ram[24454]  = 1;
  ram[24455]  = 0;
  ram[24456]  = 0;
  ram[24457]  = 1;
  ram[24458]  = 1;
  ram[24459]  = 0;
  ram[24460]  = 0;
  ram[24461]  = 1;
  ram[24462]  = 1;
  ram[24463]  = 1;
  ram[24464]  = 0;
  ram[24465]  = 0;
  ram[24466]  = 1;
  ram[24467]  = 1;
  ram[24468]  = 1;
  ram[24469]  = 1;
  ram[24470]  = 1;
  ram[24471]  = 0;
  ram[24472]  = 1;
  ram[24473]  = 1;
  ram[24474]  = 1;
  ram[24475]  = 1;
  ram[24476]  = 1;
  ram[24477]  = 1;
  ram[24478]  = 1;
  ram[24479]  = 1;
  ram[24480]  = 0;
  ram[24481]  = 0;
  ram[24482]  = 1;
  ram[24483]  = 1;
  ram[24484]  = 1;
  ram[24485]  = 1;
  ram[24486]  = 0;
  ram[24487]  = 0;
  ram[24488]  = 1;
  ram[24489]  = 1;
  ram[24490]  = 1;
  ram[24491]  = 0;
  ram[24492]  = 0;
  ram[24493]  = 1;
  ram[24494]  = 1;
  ram[24495]  = 1;
  ram[24496]  = 1;
  ram[24497]  = 1;
  ram[24498]  = 1;
  ram[24499]  = 1;
  ram[24500]  = 1;
  ram[24501]  = 0;
  ram[24502]  = 0;
  ram[24503]  = 1;
  ram[24504]  = 1;
  ram[24505]  = 1;
  ram[24506]  = 1;
  ram[24507]  = 1;
  ram[24508]  = 0;
  ram[24509]  = 0;
  ram[24510]  = 1;
  ram[24511]  = 1;
  ram[24512]  = 0;
  ram[24513]  = 0;
  ram[24514]  = 1;
  ram[24515]  = 1;
  ram[24516]  = 1;
  ram[24517]  = 0;
  ram[24518]  = 1;
  ram[24519]  = 1;
  ram[24520]  = 1;
  ram[24521]  = 0;
  ram[24522]  = 1;
  ram[24523]  = 1;
  ram[24524]  = 1;
  ram[24525]  = 0;
  ram[24526]  = 0;
  ram[24527]  = 1;
  ram[24528]  = 1;
  ram[24529]  = 1;
  ram[24530]  = 0;
  ram[24531]  = 0;
  ram[24532]  = 1;
  ram[24533]  = 1;
  ram[24534]  = 0;
  ram[24535]  = 1;
  ram[24536]  = 0;
  ram[24537]  = 1;
  ram[24538]  = 1;
  ram[24539]  = 1;
  ram[24540]  = 0;
  ram[24541]  = 1;
  ram[24542]  = 1;
  ram[24543]  = 1;
  ram[24544]  = 1;
  ram[24545]  = 1;
  ram[24546]  = 1;
  ram[24547]  = 0;
  ram[24548]  = 1;
  ram[24549]  = 1;
  ram[24550]  = 1;
  ram[24551]  = 1;
  ram[24552]  = 1;
  ram[24553]  = 1;
  ram[24554]  = 1;
  ram[24555]  = 1;
  ram[24556]  = 1;
  ram[24557]  = 1;
  ram[24558]  = 1;
  ram[24559]  = 1;
  ram[24560]  = 1;
  ram[24561]  = 1;
  ram[24562]  = 1;
  ram[24563]  = 1;
  ram[24564]  = 1;
  ram[24565]  = 1;
  ram[24566]  = 1;
  ram[24567]  = 1;
  ram[24568]  = 1;
  ram[24569]  = 1;
  ram[24570]  = 1;
  ram[24571]  = 1;
  ram[24572]  = 1;
  ram[24573]  = 1;
  ram[24574]  = 1;
  ram[24575]  = 1;
  ram[24576]  = 1;
  ram[24577]  = 1;
  ram[24578]  = 1;
  ram[24579]  = 1;
  ram[24580]  = 1;
  ram[24581]  = 1;
  ram[24582]  = 1;
  ram[24583]  = 1;
  ram[24584]  = 1;
  ram[24585]  = 1;
  ram[24586]  = 1;
  ram[24587]  = 1;
  ram[24588]  = 1;
  ram[24589]  = 1;
  ram[24590]  = 1;
  ram[24591]  = 1;
  ram[24592]  = 1;
  ram[24593]  = 1;
  ram[24594]  = 1;
  ram[24595]  = 1;
  ram[24596]  = 1;
  ram[24597]  = 1;
  ram[24598]  = 1;
  ram[24599]  = 1;
  ram[24600]  = 1;
  ram[24601]  = 1;
  ram[24602]  = 1;
  ram[24603]  = 1;
  ram[24604]  = 1;
  ram[24605]  = 1;
  ram[24606]  = 1;
  ram[24607]  = 1;
  ram[24608]  = 1;
  ram[24609]  = 1;
  ram[24610]  = 1;
  ram[24611]  = 1;
  ram[24612]  = 1;
  ram[24613]  = 1;
  ram[24614]  = 1;
  ram[24615]  = 1;
  ram[24616]  = 1;
  ram[24617]  = 1;
  ram[24618]  = 1;
  ram[24619]  = 1;
  ram[24620]  = 1;
  ram[24621]  = 1;
  ram[24622]  = 1;
  ram[24623]  = 1;
  ram[24624]  = 1;
  ram[24625]  = 1;
  ram[24626]  = 1;
  ram[24627]  = 1;
  ram[24628]  = 1;
  ram[24629]  = 1;
  ram[24630]  = 1;
  ram[24631]  = 1;
  ram[24632]  = 1;
  ram[24633]  = 1;
  ram[24634]  = 1;
  ram[24635]  = 1;
  ram[24636]  = 1;
  ram[24637]  = 1;
  ram[24638]  = 1;
  ram[24639]  = 1;
  ram[24640]  = 1;
  ram[24641]  = 1;
  ram[24642]  = 1;
  ram[24643]  = 1;
  ram[24644]  = 1;
  ram[24645]  = 0;
  ram[24646]  = 1;
  ram[24647]  = 1;
  ram[24648]  = 1;
  ram[24649]  = 1;
  ram[24650]  = 1;
  ram[24651]  = 1;
  ram[24652]  = 1;
  ram[24653]  = 1;
  ram[24654]  = 1;
  ram[24655]  = 0;
  ram[24656]  = 1;
  ram[24657]  = 1;
  ram[24658]  = 1;
  ram[24659]  = 1;
  ram[24660]  = 1;
  ram[24661]  = 1;
  ram[24662]  = 1;
  ram[24663]  = 0;
  ram[24664]  = 0;
  ram[24665]  = 0;
  ram[24666]  = 0;
  ram[24667]  = 1;
  ram[24668]  = 1;
  ram[24669]  = 1;
  ram[24670]  = 1;
  ram[24671]  = 0;
  ram[24672]  = 0;
  ram[24673]  = 0;
  ram[24674]  = 0;
  ram[24675]  = 1;
  ram[24676]  = 1;
  ram[24677]  = 1;
  ram[24678]  = 0;
  ram[24679]  = 0;
  ram[24680]  = 0;
  ram[24681]  = 0;
  ram[24682]  = 0;
  ram[24683]  = 1;
  ram[24684]  = 1;
  ram[24685]  = 1;
  ram[24686]  = 1;
  ram[24687]  = 1;
  ram[24688]  = 1;
  ram[24689]  = 1;
  ram[24690]  = 1;
  ram[24691]  = 1;
  ram[24692]  = 0;
  ram[24693]  = 0;
  ram[24694]  = 0;
  ram[24695]  = 1;
  ram[24696]  = 1;
  ram[24697]  = 0;
  ram[24698]  = 1;
  ram[24699]  = 1;
  ram[24700]  = 1;
  ram[24701]  = 1;
  ram[24702]  = 1;
  ram[24703]  = 0;
  ram[24704]  = 1;
  ram[24705]  = 1;
  ram[24706]  = 1;
  ram[24707]  = 1;
  ram[24708]  = 0;
  ram[24709]  = 0;
  ram[24710]  = 0;
  ram[24711]  = 0;
  ram[24712]  = 0;
  ram[24713]  = 1;
  ram[24714]  = 1;
  ram[24715]  = 1;
  ram[24716]  = 1;
  ram[24717]  = 1;
  ram[24718]  = 1;
  ram[24719]  = 1;
  ram[24720]  = 1;
  ram[24721]  = 1;
  ram[24722]  = 0;
  ram[24723]  = 0;
  ram[24724]  = 0;
  ram[24725]  = 0;
  ram[24726]  = 0;
  ram[24727]  = 1;
  ram[24728]  = 1;
  ram[24729]  = 1;
  ram[24730]  = 1;
  ram[24731]  = 1;
  ram[24732]  = 1;
  ram[24733]  = 0;
  ram[24734]  = 0;
  ram[24735]  = 0;
  ram[24736]  = 0;
  ram[24737]  = 1;
  ram[24738]  = 0;
  ram[24739]  = 1;
  ram[24740]  = 1;
  ram[24741]  = 1;
  ram[24742]  = 1;
  ram[24743]  = 0;
  ram[24744]  = 0;
  ram[24745]  = 0;
  ram[24746]  = 1;
  ram[24747]  = 1;
  ram[24748]  = 1;
  ram[24749]  = 0;
  ram[24750]  = 0;
  ram[24751]  = 0;
  ram[24752]  = 1;
  ram[24753]  = 1;
  ram[24754]  = 1;
  ram[24755]  = 0;
  ram[24756]  = 0;
  ram[24757]  = 0;
  ram[24758]  = 0;
  ram[24759]  = 0;
  ram[24760]  = 1;
  ram[24761]  = 1;
  ram[24762]  = 1;
  ram[24763]  = 1;
  ram[24764]  = 0;
  ram[24765]  = 0;
  ram[24766]  = 1;
  ram[24767]  = 1;
  ram[24768]  = 1;
  ram[24769]  = 1;
  ram[24770]  = 1;
  ram[24771]  = 0;
  ram[24772]  = 1;
  ram[24773]  = 1;
  ram[24774]  = 1;
  ram[24775]  = 1;
  ram[24776]  = 1;
  ram[24777]  = 1;
  ram[24778]  = 1;
  ram[24779]  = 1;
  ram[24780]  = 1;
  ram[24781]  = 0;
  ram[24782]  = 0;
  ram[24783]  = 0;
  ram[24784]  = 1;
  ram[24785]  = 1;
  ram[24786]  = 1;
  ram[24787]  = 0;
  ram[24788]  = 0;
  ram[24789]  = 0;
  ram[24790]  = 0;
  ram[24791]  = 0;
  ram[24792]  = 1;
  ram[24793]  = 1;
  ram[24794]  = 1;
  ram[24795]  = 1;
  ram[24796]  = 1;
  ram[24797]  = 1;
  ram[24798]  = 1;
  ram[24799]  = 1;
  ram[24800]  = 1;
  ram[24801]  = 0;
  ram[24802]  = 0;
  ram[24803]  = 1;
  ram[24804]  = 1;
  ram[24805]  = 1;
  ram[24806]  = 1;
  ram[24807]  = 1;
  ram[24808]  = 1;
  ram[24809]  = 0;
  ram[24810]  = 0;
  ram[24811]  = 0;
  ram[24812]  = 0;
  ram[24813]  = 1;
  ram[24814]  = 1;
  ram[24815]  = 1;
  ram[24816]  = 1;
  ram[24817]  = 0;
  ram[24818]  = 0;
  ram[24819]  = 0;
  ram[24820]  = 0;
  ram[24821]  = 0;
  ram[24822]  = 1;
  ram[24823]  = 1;
  ram[24824]  = 1;
  ram[24825]  = 1;
  ram[24826]  = 0;
  ram[24827]  = 0;
  ram[24828]  = 0;
  ram[24829]  = 1;
  ram[24830]  = 1;
  ram[24831]  = 0;
  ram[24832]  = 0;
  ram[24833]  = 0;
  ram[24834]  = 0;
  ram[24835]  = 1;
  ram[24836]  = 0;
  ram[24837]  = 1;
  ram[24838]  = 1;
  ram[24839]  = 1;
  ram[24840]  = 0;
  ram[24841]  = 1;
  ram[24842]  = 1;
  ram[24843]  = 1;
  ram[24844]  = 1;
  ram[24845]  = 1;
  ram[24846]  = 1;
  ram[24847]  = 0;
  ram[24848]  = 0;
  ram[24849]  = 0;
  ram[24850]  = 1;
  ram[24851]  = 1;
  ram[24852]  = 1;
  ram[24853]  = 1;
  ram[24854]  = 1;
  ram[24855]  = 1;
  ram[24856]  = 1;
  ram[24857]  = 1;
  ram[24858]  = 1;
  ram[24859]  = 1;
  ram[24860]  = 1;
  ram[24861]  = 1;
  ram[24862]  = 1;
  ram[24863]  = 1;
  ram[24864]  = 1;
  ram[24865]  = 1;
  ram[24866]  = 1;
  ram[24867]  = 1;
  ram[24868]  = 1;
  ram[24869]  = 1;
  ram[24870]  = 1;
  ram[24871]  = 1;
  ram[24872]  = 1;
  ram[24873]  = 1;
  ram[24874]  = 1;
  ram[24875]  = 1;
  ram[24876]  = 1;
  ram[24877]  = 1;
  ram[24878]  = 1;
  ram[24879]  = 1;
  ram[24880]  = 1;
  ram[24881]  = 1;
  ram[24882]  = 1;
  ram[24883]  = 1;
  ram[24884]  = 1;
  ram[24885]  = 1;
  ram[24886]  = 1;
  ram[24887]  = 1;
  ram[24888]  = 1;
  ram[24889]  = 1;
  ram[24890]  = 1;
  ram[24891]  = 1;
  ram[24892]  = 1;
  ram[24893]  = 1;
  ram[24894]  = 1;
  ram[24895]  = 1;
  ram[24896]  = 1;
  ram[24897]  = 1;
  ram[24898]  = 1;
  ram[24899]  = 1;
  ram[24900]  = 1;
  ram[24901]  = 1;
  ram[24902]  = 1;
  ram[24903]  = 1;
  ram[24904]  = 1;
  ram[24905]  = 1;
  ram[24906]  = 1;
  ram[24907]  = 1;
  ram[24908]  = 1;
  ram[24909]  = 1;
  ram[24910]  = 1;
  ram[24911]  = 1;
  ram[24912]  = 1;
  ram[24913]  = 1;
  ram[24914]  = 1;
  ram[24915]  = 1;
  ram[24916]  = 1;
  ram[24917]  = 1;
  ram[24918]  = 1;
  ram[24919]  = 1;
  ram[24920]  = 1;
  ram[24921]  = 1;
  ram[24922]  = 1;
  ram[24923]  = 1;
  ram[24924]  = 1;
  ram[24925]  = 1;
  ram[24926]  = 1;
  ram[24927]  = 1;
  ram[24928]  = 1;
  ram[24929]  = 1;
  ram[24930]  = 1;
  ram[24931]  = 1;
  ram[24932]  = 1;
  ram[24933]  = 1;
  ram[24934]  = 1;
  ram[24935]  = 1;
  ram[24936]  = 1;
  ram[24937]  = 1;
  ram[24938]  = 1;
  ram[24939]  = 1;
  ram[24940]  = 1;
  ram[24941]  = 1;
  ram[24942]  = 1;
  ram[24943]  = 1;
  ram[24944]  = 1;
  ram[24945]  = 1;
  ram[24946]  = 1;
  ram[24947]  = 1;
  ram[24948]  = 1;
  ram[24949]  = 1;
  ram[24950]  = 1;
  ram[24951]  = 1;
  ram[24952]  = 1;
  ram[24953]  = 1;
  ram[24954]  = 1;
  ram[24955]  = 1;
  ram[24956]  = 1;
  ram[24957]  = 1;
  ram[24958]  = 1;
  ram[24959]  = 1;
  ram[24960]  = 1;
  ram[24961]  = 1;
  ram[24962]  = 1;
  ram[24963]  = 1;
  ram[24964]  = 1;
  ram[24965]  = 1;
  ram[24966]  = 1;
  ram[24967]  = 1;
  ram[24968]  = 1;
  ram[24969]  = 1;
  ram[24970]  = 1;
  ram[24971]  = 1;
  ram[24972]  = 1;
  ram[24973]  = 1;
  ram[24974]  = 1;
  ram[24975]  = 1;
  ram[24976]  = 1;
  ram[24977]  = 1;
  ram[24978]  = 1;
  ram[24979]  = 1;
  ram[24980]  = 1;
  ram[24981]  = 1;
  ram[24982]  = 1;
  ram[24983]  = 1;
  ram[24984]  = 1;
  ram[24985]  = 1;
  ram[24986]  = 1;
  ram[24987]  = 1;
  ram[24988]  = 1;
  ram[24989]  = 1;
  ram[24990]  = 1;
  ram[24991]  = 1;
  ram[24992]  = 1;
  ram[24993]  = 1;
  ram[24994]  = 1;
  ram[24995]  = 1;
  ram[24996]  = 1;
  ram[24997]  = 1;
  ram[24998]  = 1;
  ram[24999]  = 1;
  ram[25000]  = 1;
  ram[25001]  = 1;
  ram[25002]  = 1;
  ram[25003]  = 1;
  ram[25004]  = 1;
  ram[25005]  = 1;
  ram[25006]  = 1;
  ram[25007]  = 1;
  ram[25008]  = 1;
  ram[25009]  = 1;
  ram[25010]  = 1;
  ram[25011]  = 1;
  ram[25012]  = 1;
  ram[25013]  = 1;
  ram[25014]  = 1;
  ram[25015]  = 1;
  ram[25016]  = 1;
  ram[25017]  = 1;
  ram[25018]  = 1;
  ram[25019]  = 1;
  ram[25020]  = 1;
  ram[25021]  = 1;
  ram[25022]  = 1;
  ram[25023]  = 1;
  ram[25024]  = 1;
  ram[25025]  = 1;
  ram[25026]  = 1;
  ram[25027]  = 1;
  ram[25028]  = 1;
  ram[25029]  = 1;
  ram[25030]  = 1;
  ram[25031]  = 1;
  ram[25032]  = 1;
  ram[25033]  = 1;
  ram[25034]  = 1;
  ram[25035]  = 1;
  ram[25036]  = 1;
  ram[25037]  = 1;
  ram[25038]  = 1;
  ram[25039]  = 1;
  ram[25040]  = 1;
  ram[25041]  = 1;
  ram[25042]  = 1;
  ram[25043]  = 1;
  ram[25044]  = 1;
  ram[25045]  = 1;
  ram[25046]  = 1;
  ram[25047]  = 1;
  ram[25048]  = 1;
  ram[25049]  = 1;
  ram[25050]  = 1;
  ram[25051]  = 1;
  ram[25052]  = 1;
  ram[25053]  = 1;
  ram[25054]  = 1;
  ram[25055]  = 1;
  ram[25056]  = 1;
  ram[25057]  = 1;
  ram[25058]  = 1;
  ram[25059]  = 1;
  ram[25060]  = 1;
  ram[25061]  = 1;
  ram[25062]  = 1;
  ram[25063]  = 1;
  ram[25064]  = 1;
  ram[25065]  = 1;
  ram[25066]  = 1;
  ram[25067]  = 1;
  ram[25068]  = 1;
  ram[25069]  = 1;
  ram[25070]  = 1;
  ram[25071]  = 1;
  ram[25072]  = 1;
  ram[25073]  = 1;
  ram[25074]  = 1;
  ram[25075]  = 1;
  ram[25076]  = 1;
  ram[25077]  = 1;
  ram[25078]  = 1;
  ram[25079]  = 1;
  ram[25080]  = 1;
  ram[25081]  = 1;
  ram[25082]  = 1;
  ram[25083]  = 1;
  ram[25084]  = 1;
  ram[25085]  = 1;
  ram[25086]  = 1;
  ram[25087]  = 1;
  ram[25088]  = 1;
  ram[25089]  = 1;
  ram[25090]  = 1;
  ram[25091]  = 1;
  ram[25092]  = 1;
  ram[25093]  = 1;
  ram[25094]  = 1;
  ram[25095]  = 1;
  ram[25096]  = 1;
  ram[25097]  = 1;
  ram[25098]  = 1;
  ram[25099]  = 1;
  ram[25100]  = 1;
  ram[25101]  = 1;
  ram[25102]  = 1;
  ram[25103]  = 1;
  ram[25104]  = 1;
  ram[25105]  = 1;
  ram[25106]  = 1;
  ram[25107]  = 1;
  ram[25108]  = 1;
  ram[25109]  = 1;
  ram[25110]  = 1;
  ram[25111]  = 1;
  ram[25112]  = 1;
  ram[25113]  = 1;
  ram[25114]  = 1;
  ram[25115]  = 1;
  ram[25116]  = 1;
  ram[25117]  = 1;
  ram[25118]  = 1;
  ram[25119]  = 1;
  ram[25120]  = 1;
  ram[25121]  = 1;
  ram[25122]  = 1;
  ram[25123]  = 1;
  ram[25124]  = 1;
  ram[25125]  = 1;
  ram[25126]  = 1;
  ram[25127]  = 1;
  ram[25128]  = 1;
  ram[25129]  = 1;
  ram[25130]  = 1;
  ram[25131]  = 1;
  ram[25132]  = 1;
  ram[25133]  = 1;
  ram[25134]  = 1;
  ram[25135]  = 1;
  ram[25136]  = 1;
  ram[25137]  = 1;
  ram[25138]  = 1;
  ram[25139]  = 1;
  ram[25140]  = 1;
  ram[25141]  = 1;
  ram[25142]  = 1;
  ram[25143]  = 1;
  ram[25144]  = 1;
  ram[25145]  = 1;
  ram[25146]  = 1;
  ram[25147]  = 1;
  ram[25148]  = 1;
  ram[25149]  = 1;
  ram[25150]  = 1;
  ram[25151]  = 1;
  ram[25152]  = 1;
  ram[25153]  = 1;
  ram[25154]  = 1;
  ram[25155]  = 1;
  ram[25156]  = 1;
  ram[25157]  = 1;
  ram[25158]  = 1;
  ram[25159]  = 1;
  ram[25160]  = 1;
  ram[25161]  = 1;
  ram[25162]  = 1;
  ram[25163]  = 1;
  ram[25164]  = 1;
  ram[25165]  = 1;
  ram[25166]  = 1;
  ram[25167]  = 1;
  ram[25168]  = 1;
  ram[25169]  = 1;
  ram[25170]  = 1;
  ram[25171]  = 1;
  ram[25172]  = 1;
  ram[25173]  = 1;
  ram[25174]  = 1;
  ram[25175]  = 1;
  ram[25176]  = 1;
  ram[25177]  = 1;
  ram[25178]  = 1;
  ram[25179]  = 1;
  ram[25180]  = 1;
  ram[25181]  = 1;
  ram[25182]  = 1;
  ram[25183]  = 1;
  ram[25184]  = 1;
  ram[25185]  = 1;
  ram[25186]  = 1;
  ram[25187]  = 1;
  ram[25188]  = 1;
  ram[25189]  = 1;
  ram[25190]  = 1;
  ram[25191]  = 1;
  ram[25192]  = 1;
  ram[25193]  = 1;
  ram[25194]  = 1;
  ram[25195]  = 1;
  ram[25196]  = 1;
  ram[25197]  = 1;
  ram[25198]  = 1;
  ram[25199]  = 1;
  ram[25200]  = 1;
  ram[25201]  = 1;
  ram[25202]  = 1;
  ram[25203]  = 1;
  ram[25204]  = 1;
  ram[25205]  = 1;
  ram[25206]  = 1;
  ram[25207]  = 1;
  ram[25208]  = 1;
  ram[25209]  = 1;
  ram[25210]  = 1;
  ram[25211]  = 1;
  ram[25212]  = 1;
  ram[25213]  = 1;
  ram[25214]  = 1;
  ram[25215]  = 1;
  ram[25216]  = 1;
  ram[25217]  = 1;
  ram[25218]  = 1;
  ram[25219]  = 1;
  ram[25220]  = 1;
  ram[25221]  = 1;
  ram[25222]  = 1;
  ram[25223]  = 1;
  ram[25224]  = 1;
  ram[25225]  = 1;
  ram[25226]  = 1;
  ram[25227]  = 1;
  ram[25228]  = 1;
  ram[25229]  = 1;
  ram[25230]  = 1;
  ram[25231]  = 1;
  ram[25232]  = 1;
  ram[25233]  = 1;
  ram[25234]  = 1;
  ram[25235]  = 1;
  ram[25236]  = 1;
  ram[25237]  = 1;
  ram[25238]  = 1;
  ram[25239]  = 1;
  ram[25240]  = 1;
  ram[25241]  = 1;
  ram[25242]  = 1;
  ram[25243]  = 1;
  ram[25244]  = 1;
  ram[25245]  = 1;
  ram[25246]  = 1;
  ram[25247]  = 1;
  ram[25248]  = 1;
  ram[25249]  = 1;
  ram[25250]  = 1;
  ram[25251]  = 1;
  ram[25252]  = 1;
  ram[25253]  = 1;
  ram[25254]  = 1;
  ram[25255]  = 1;
  ram[25256]  = 1;
  ram[25257]  = 1;
  ram[25258]  = 1;
  ram[25259]  = 1;
  ram[25260]  = 1;
  ram[25261]  = 1;
  ram[25262]  = 1;
  ram[25263]  = 1;
  ram[25264]  = 1;
  ram[25265]  = 1;
  ram[25266]  = 1;
  ram[25267]  = 1;
  ram[25268]  = 1;
  ram[25269]  = 1;
  ram[25270]  = 1;
  ram[25271]  = 1;
  ram[25272]  = 1;
  ram[25273]  = 1;
  ram[25274]  = 1;
  ram[25275]  = 1;
  ram[25276]  = 1;
  ram[25277]  = 1;
  ram[25278]  = 1;
  ram[25279]  = 1;
  ram[25280]  = 1;
  ram[25281]  = 1;
  ram[25282]  = 1;
  ram[25283]  = 1;
  ram[25284]  = 1;
  ram[25285]  = 1;
  ram[25286]  = 1;
  ram[25287]  = 1;
  ram[25288]  = 1;
  ram[25289]  = 1;
  ram[25290]  = 1;
  ram[25291]  = 1;
  ram[25292]  = 1;
  ram[25293]  = 1;
  ram[25294]  = 1;
  ram[25295]  = 1;
  ram[25296]  = 1;
  ram[25297]  = 1;
  ram[25298]  = 1;
  ram[25299]  = 1;
  ram[25300]  = 1;
  ram[25301]  = 1;
  ram[25302]  = 1;
  ram[25303]  = 1;
  ram[25304]  = 1;
  ram[25305]  = 1;
  ram[25306]  = 1;
  ram[25307]  = 1;
  ram[25308]  = 1;
  ram[25309]  = 1;
  ram[25310]  = 1;
  ram[25311]  = 1;
  ram[25312]  = 1;
  ram[25313]  = 1;
  ram[25314]  = 1;
  ram[25315]  = 1;
  ram[25316]  = 1;
  ram[25317]  = 1;
  ram[25318]  = 1;
  ram[25319]  = 1;
  ram[25320]  = 1;
  ram[25321]  = 1;
  ram[25322]  = 1;
  ram[25323]  = 1;
  ram[25324]  = 1;
  ram[25325]  = 1;
  ram[25326]  = 1;
  ram[25327]  = 1;
  ram[25328]  = 1;
  ram[25329]  = 1;
  ram[25330]  = 1;
  ram[25331]  = 1;
  ram[25332]  = 1;
  ram[25333]  = 1;
  ram[25334]  = 1;
  ram[25335]  = 1;
  ram[25336]  = 1;
  ram[25337]  = 1;
  ram[25338]  = 1;
  ram[25339]  = 1;
  ram[25340]  = 1;
  ram[25341]  = 1;
  ram[25342]  = 1;
  ram[25343]  = 1;
  ram[25344]  = 1;
  ram[25345]  = 1;
  ram[25346]  = 1;
  ram[25347]  = 1;
  ram[25348]  = 1;
  ram[25349]  = 1;
  ram[25350]  = 1;
  ram[25351]  = 1;
  ram[25352]  = 1;
  ram[25353]  = 1;
  ram[25354]  = 1;
  ram[25355]  = 1;
  ram[25356]  = 1;
  ram[25357]  = 1;
  ram[25358]  = 1;
  ram[25359]  = 1;
  ram[25360]  = 1;
  ram[25361]  = 1;
  ram[25362]  = 1;
  ram[25363]  = 1;
  ram[25364]  = 1;
  ram[25365]  = 1;
  ram[25366]  = 1;
  ram[25367]  = 1;
  ram[25368]  = 1;
  ram[25369]  = 1;
  ram[25370]  = 1;
  ram[25371]  = 1;
  ram[25372]  = 1;
  ram[25373]  = 1;
  ram[25374]  = 1;
  ram[25375]  = 1;
  ram[25376]  = 1;
  ram[25377]  = 1;
  ram[25378]  = 1;
  ram[25379]  = 1;
  ram[25380]  = 1;
  ram[25381]  = 1;
  ram[25382]  = 1;
  ram[25383]  = 1;
  ram[25384]  = 1;
  ram[25385]  = 1;
  ram[25386]  = 1;
  ram[25387]  = 1;
  ram[25388]  = 1;
  ram[25389]  = 1;
  ram[25390]  = 1;
  ram[25391]  = 1;
  ram[25392]  = 1;
  ram[25393]  = 1;
  ram[25394]  = 1;
  ram[25395]  = 1;
  ram[25396]  = 1;
  ram[25397]  = 1;
  ram[25398]  = 1;
  ram[25399]  = 1;
  ram[25400]  = 1;
  ram[25401]  = 1;
  ram[25402]  = 1;
  ram[25403]  = 1;
  ram[25404]  = 1;
  ram[25405]  = 1;
  ram[25406]  = 1;
  ram[25407]  = 1;
  ram[25408]  = 1;
  ram[25409]  = 1;
  ram[25410]  = 1;
  ram[25411]  = 1;
  ram[25412]  = 1;
  ram[25413]  = 1;
  ram[25414]  = 1;
  ram[25415]  = 1;
  ram[25416]  = 1;
  ram[25417]  = 1;
  ram[25418]  = 1;
  ram[25419]  = 1;
  ram[25420]  = 1;
  ram[25421]  = 1;
  ram[25422]  = 1;
  ram[25423]  = 1;
  ram[25424]  = 1;
  ram[25425]  = 1;
  ram[25426]  = 1;
  ram[25427]  = 1;
  ram[25428]  = 1;
  ram[25429]  = 1;
  ram[25430]  = 1;
  ram[25431]  = 1;
  ram[25432]  = 1;
  ram[25433]  = 1;
  ram[25434]  = 1;
  ram[25435]  = 1;
  ram[25436]  = 1;
  ram[25437]  = 1;
  ram[25438]  = 1;
  ram[25439]  = 1;
  ram[25440]  = 1;
  ram[25441]  = 1;
  ram[25442]  = 1;
  ram[25443]  = 1;
  ram[25444]  = 1;
  ram[25445]  = 1;
  ram[25446]  = 1;
  ram[25447]  = 1;
  ram[25448]  = 1;
  ram[25449]  = 1;
  ram[25450]  = 1;
  ram[25451]  = 1;
  ram[25452]  = 1;
  ram[25453]  = 1;
  ram[25454]  = 1;
  ram[25455]  = 1;
  ram[25456]  = 1;
  ram[25457]  = 1;
  ram[25458]  = 1;
  ram[25459]  = 1;
  ram[25460]  = 1;
  ram[25461]  = 1;
  ram[25462]  = 1;
  ram[25463]  = 1;
  ram[25464]  = 1;
  ram[25465]  = 1;
  ram[25466]  = 1;
  ram[25467]  = 1;
  ram[25468]  = 1;
  ram[25469]  = 1;
  ram[25470]  = 1;
  ram[25471]  = 1;
  ram[25472]  = 1;
  ram[25473]  = 1;
  ram[25474]  = 1;
  ram[25475]  = 1;
  ram[25476]  = 1;
  ram[25477]  = 1;
  ram[25478]  = 1;
  ram[25479]  = 1;
  ram[25480]  = 1;
  ram[25481]  = 1;
  ram[25482]  = 1;
  ram[25483]  = 1;
  ram[25484]  = 1;
  ram[25485]  = 1;
  ram[25486]  = 1;
  ram[25487]  = 1;
  ram[25488]  = 1;
  ram[25489]  = 1;
  ram[25490]  = 1;
  ram[25491]  = 1;
  ram[25492]  = 1;
  ram[25493]  = 1;
  ram[25494]  = 1;
  ram[25495]  = 1;
  ram[25496]  = 1;
  ram[25497]  = 1;
  ram[25498]  = 1;
  ram[25499]  = 1;
  ram[25500]  = 1;
  ram[25501]  = 1;
  ram[25502]  = 1;
  ram[25503]  = 1;
  ram[25504]  = 1;
  ram[25505]  = 1;
  ram[25506]  = 1;
  ram[25507]  = 1;
  ram[25508]  = 1;
  ram[25509]  = 1;
  ram[25510]  = 1;
  ram[25511]  = 1;
  ram[25512]  = 1;
  ram[25513]  = 1;
  ram[25514]  = 1;
  ram[25515]  = 1;
  ram[25516]  = 1;
  ram[25517]  = 1;
  ram[25518]  = 1;
  ram[25519]  = 1;
  ram[25520]  = 1;
  ram[25521]  = 1;
  ram[25522]  = 1;
  ram[25523]  = 1;
  ram[25524]  = 1;
  ram[25525]  = 1;
  ram[25526]  = 1;
  ram[25527]  = 1;
  ram[25528]  = 1;
  ram[25529]  = 1;
  ram[25530]  = 1;
  ram[25531]  = 1;
  ram[25532]  = 1;
  ram[25533]  = 1;
  ram[25534]  = 1;
  ram[25535]  = 1;
  ram[25536]  = 1;
  ram[25537]  = 1;
  ram[25538]  = 1;
  ram[25539]  = 1;
  ram[25540]  = 1;
  ram[25541]  = 1;
  ram[25542]  = 1;
  ram[25543]  = 1;
  ram[25544]  = 1;
  ram[25545]  = 1;
  ram[25546]  = 1;
  ram[25547]  = 1;
  ram[25548]  = 1;
  ram[25549]  = 1;
  ram[25550]  = 1;
  ram[25551]  = 1;
  ram[25552]  = 1;
  ram[25553]  = 1;
  ram[25554]  = 1;
  ram[25555]  = 1;
  ram[25556]  = 1;
  ram[25557]  = 1;
  ram[25558]  = 1;
  ram[25559]  = 1;
  ram[25560]  = 1;
  ram[25561]  = 1;
  ram[25562]  = 1;
  ram[25563]  = 1;
  ram[25564]  = 1;
  ram[25565]  = 1;
  ram[25566]  = 1;
  ram[25567]  = 1;
  ram[25568]  = 1;
  ram[25569]  = 1;
  ram[25570]  = 1;
  ram[25571]  = 1;
  ram[25572]  = 1;
  ram[25573]  = 1;
  ram[25574]  = 1;
  ram[25575]  = 1;
  ram[25576]  = 1;
  ram[25577]  = 1;
  ram[25578]  = 1;
  ram[25579]  = 1;
  ram[25580]  = 1;
  ram[25581]  = 1;
  ram[25582]  = 1;
  ram[25583]  = 1;
  ram[25584]  = 1;
  ram[25585]  = 1;
  ram[25586]  = 1;
  ram[25587]  = 1;
  ram[25588]  = 1;
  ram[25589]  = 1;
  ram[25590]  = 1;
  ram[25591]  = 1;
  ram[25592]  = 1;
  ram[25593]  = 1;
  ram[25594]  = 1;
  ram[25595]  = 1;
  ram[25596]  = 1;
  ram[25597]  = 1;
  ram[25598]  = 1;
  ram[25599]  = 1;
  ram[25600]  = 1;
  ram[25601]  = 1;
  ram[25602]  = 1;
  ram[25603]  = 1;
  ram[25604]  = 1;
  ram[25605]  = 1;
  ram[25606]  = 1;
  ram[25607]  = 1;
  ram[25608]  = 1;
  ram[25609]  = 1;
  ram[25610]  = 1;
  ram[25611]  = 1;
  ram[25612]  = 1;
  ram[25613]  = 1;
  ram[25614]  = 1;
  ram[25615]  = 1;
  ram[25616]  = 1;
  ram[25617]  = 1;
  ram[25618]  = 1;
  ram[25619]  = 1;
  ram[25620]  = 1;
  ram[25621]  = 1;
  ram[25622]  = 1;
  ram[25623]  = 1;
  ram[25624]  = 1;
  ram[25625]  = 1;
  ram[25626]  = 1;
  ram[25627]  = 1;
  ram[25628]  = 1;
  ram[25629]  = 1;
  ram[25630]  = 1;
  ram[25631]  = 1;
  ram[25632]  = 1;
  ram[25633]  = 1;
  ram[25634]  = 1;
  ram[25635]  = 1;
  ram[25636]  = 1;
  ram[25637]  = 1;
  ram[25638]  = 1;
  ram[25639]  = 1;
  ram[25640]  = 1;
  ram[25641]  = 1;
  ram[25642]  = 1;
  ram[25643]  = 1;
  ram[25644]  = 1;
  ram[25645]  = 1;
  ram[25646]  = 1;
  ram[25647]  = 1;
  ram[25648]  = 1;
  ram[25649]  = 1;
  ram[25650]  = 1;
  ram[25651]  = 1;
  ram[25652]  = 1;
  ram[25653]  = 1;
  ram[25654]  = 1;
  ram[25655]  = 1;
  ram[25656]  = 1;
  ram[25657]  = 1;
  ram[25658]  = 1;
  ram[25659]  = 1;
  ram[25660]  = 1;
  ram[25661]  = 1;
  ram[25662]  = 1;
  ram[25663]  = 1;
  ram[25664]  = 1;
  ram[25665]  = 1;
  ram[25666]  = 1;
  ram[25667]  = 1;
  ram[25668]  = 1;
  ram[25669]  = 1;
  ram[25670]  = 1;
  ram[25671]  = 1;
  ram[25672]  = 1;
  ram[25673]  = 1;
  ram[25674]  = 1;
  ram[25675]  = 1;
  ram[25676]  = 1;
  ram[25677]  = 1;
  ram[25678]  = 1;
  ram[25679]  = 1;
  ram[25680]  = 1;
  ram[25681]  = 1;
  ram[25682]  = 1;
  ram[25683]  = 1;
  ram[25684]  = 1;
  ram[25685]  = 1;
  ram[25686]  = 1;
  ram[25687]  = 1;
  ram[25688]  = 1;
  ram[25689]  = 1;
  ram[25690]  = 1;
  ram[25691]  = 1;
  ram[25692]  = 1;
  ram[25693]  = 1;
  ram[25694]  = 1;
  ram[25695]  = 1;
  ram[25696]  = 1;
  ram[25697]  = 1;
  ram[25698]  = 1;
  ram[25699]  = 1;
  ram[25700]  = 1;
  ram[25701]  = 1;
  ram[25702]  = 1;
  ram[25703]  = 1;
  ram[25704]  = 1;
  ram[25705]  = 1;
  ram[25706]  = 1;
  ram[25707]  = 1;
  ram[25708]  = 1;
  ram[25709]  = 1;
  ram[25710]  = 1;
  ram[25711]  = 1;
  ram[25712]  = 1;
  ram[25713]  = 1;
  ram[25714]  = 1;
  ram[25715]  = 1;
  ram[25716]  = 1;
  ram[25717]  = 1;
  ram[25718]  = 1;
  ram[25719]  = 1;
  ram[25720]  = 1;
  ram[25721]  = 1;
  ram[25722]  = 1;
  ram[25723]  = 1;
  ram[25724]  = 1;
  ram[25725]  = 1;
  ram[25726]  = 1;
  ram[25727]  = 1;
  ram[25728]  = 1;
  ram[25729]  = 1;
  ram[25730]  = 1;
  ram[25731]  = 1;
  ram[25732]  = 1;
  ram[25733]  = 1;
  ram[25734]  = 1;
  ram[25735]  = 1;
  ram[25736]  = 1;
  ram[25737]  = 1;
  ram[25738]  = 1;
  ram[25739]  = 1;
  ram[25740]  = 1;
  ram[25741]  = 1;
  ram[25742]  = 1;
  ram[25743]  = 1;
  ram[25744]  = 1;
  ram[25745]  = 1;
  ram[25746]  = 1;
  ram[25747]  = 1;
  ram[25748]  = 1;
  ram[25749]  = 1;
  ram[25750]  = 1;
  ram[25751]  = 1;
  ram[25752]  = 1;
  ram[25753]  = 1;
  ram[25754]  = 1;
  ram[25755]  = 1;
  ram[25756]  = 1;
  ram[25757]  = 1;
  ram[25758]  = 1;
  ram[25759]  = 1;
  ram[25760]  = 1;
  ram[25761]  = 1;
  ram[25762]  = 1;
  ram[25763]  = 1;
  ram[25764]  = 1;
  ram[25765]  = 1;
  ram[25766]  = 1;
  ram[25767]  = 1;
  ram[25768]  = 1;
  ram[25769]  = 1;
  ram[25770]  = 1;
  ram[25771]  = 1;
  ram[25772]  = 1;
  ram[25773]  = 1;
  ram[25774]  = 1;
  ram[25775]  = 1;
  ram[25776]  = 1;
  ram[25777]  = 1;
  ram[25778]  = 1;
  ram[25779]  = 1;
  ram[25780]  = 1;
  ram[25781]  = 1;
  ram[25782]  = 1;
  ram[25783]  = 1;
  ram[25784]  = 1;
  ram[25785]  = 1;
  ram[25786]  = 1;
  ram[25787]  = 1;
  ram[25788]  = 1;
  ram[25789]  = 1;
  ram[25790]  = 1;
  ram[25791]  = 1;
  ram[25792]  = 1;
  ram[25793]  = 1;
  ram[25794]  = 1;
  ram[25795]  = 1;
  ram[25796]  = 1;
  ram[25797]  = 1;
  ram[25798]  = 1;
  ram[25799]  = 1;
  ram[25800]  = 1;
  ram[25801]  = 1;
  ram[25802]  = 1;
  ram[25803]  = 1;
  ram[25804]  = 1;
  ram[25805]  = 1;
  ram[25806]  = 1;
  ram[25807]  = 1;
  ram[25808]  = 1;
  ram[25809]  = 1;
  ram[25810]  = 1;
  ram[25811]  = 1;
  ram[25812]  = 1;
  ram[25813]  = 1;
  ram[25814]  = 1;
  ram[25815]  = 1;
  ram[25816]  = 1;
  ram[25817]  = 1;
  ram[25818]  = 1;
  ram[25819]  = 1;
  ram[25820]  = 1;
  ram[25821]  = 1;
  ram[25822]  = 1;
  ram[25823]  = 1;
  ram[25824]  = 1;
  ram[25825]  = 1;
  ram[25826]  = 1;
  ram[25827]  = 1;
  ram[25828]  = 1;
  ram[25829]  = 1;
  ram[25830]  = 1;
  ram[25831]  = 1;
  ram[25832]  = 1;
  ram[25833]  = 1;
  ram[25834]  = 1;
  ram[25835]  = 1;
  ram[25836]  = 1;
  ram[25837]  = 1;
  ram[25838]  = 1;
  ram[25839]  = 1;
  ram[25840]  = 1;
  ram[25841]  = 1;
  ram[25842]  = 1;
  ram[25843]  = 1;
  ram[25844]  = 1;
  ram[25845]  = 1;
  ram[25846]  = 1;
  ram[25847]  = 1;
  ram[25848]  = 1;
  ram[25849]  = 1;
  ram[25850]  = 1;
  ram[25851]  = 1;
  ram[25852]  = 1;
  ram[25853]  = 1;
  ram[25854]  = 1;
  ram[25855]  = 1;
  ram[25856]  = 1;
  ram[25857]  = 1;
  ram[25858]  = 1;
  ram[25859]  = 1;
  ram[25860]  = 1;
  ram[25861]  = 1;
  ram[25862]  = 1;
  ram[25863]  = 1;
  ram[25864]  = 1;
  ram[25865]  = 1;
  ram[25866]  = 1;
  ram[25867]  = 1;
  ram[25868]  = 1;
  ram[25869]  = 1;
  ram[25870]  = 1;
  ram[25871]  = 1;
  ram[25872]  = 1;
  ram[25873]  = 1;
  ram[25874]  = 1;
  ram[25875]  = 1;
  ram[25876]  = 1;
  ram[25877]  = 1;
  ram[25878]  = 1;
  ram[25879]  = 1;
  ram[25880]  = 1;
  ram[25881]  = 1;
  ram[25882]  = 1;
  ram[25883]  = 1;
  ram[25884]  = 1;
  ram[25885]  = 1;
  ram[25886]  = 1;
  ram[25887]  = 1;
  ram[25888]  = 1;
  ram[25889]  = 1;
  ram[25890]  = 1;
  ram[25891]  = 1;
  ram[25892]  = 1;
  ram[25893]  = 1;
  ram[25894]  = 1;
  ram[25895]  = 1;
  ram[25896]  = 1;
  ram[25897]  = 1;
  ram[25898]  = 1;
  ram[25899]  = 1;
  ram[25900]  = 1;
  ram[25901]  = 1;
  ram[25902]  = 1;
  ram[25903]  = 1;
  ram[25904]  = 1;
  ram[25905]  = 1;
  ram[25906]  = 1;
  ram[25907]  = 1;
  ram[25908]  = 1;
  ram[25909]  = 1;
  ram[25910]  = 1;
  ram[25911]  = 1;
  ram[25912]  = 1;
  ram[25913]  = 1;
  ram[25914]  = 1;
  ram[25915]  = 1;
  ram[25916]  = 1;
  ram[25917]  = 1;
  ram[25918]  = 1;
  ram[25919]  = 1;
  ram[25920]  = 1;
  ram[25921]  = 1;
  ram[25922]  = 1;
  ram[25923]  = 1;
  ram[25924]  = 1;
  ram[25925]  = 1;
  ram[25926]  = 1;
  ram[25927]  = 1;
  ram[25928]  = 1;
  ram[25929]  = 1;
  ram[25930]  = 1;
  ram[25931]  = 1;
  ram[25932]  = 1;
  ram[25933]  = 1;
  ram[25934]  = 1;
  ram[25935]  = 1;
  ram[25936]  = 1;
  ram[25937]  = 1;
  ram[25938]  = 1;
  ram[25939]  = 1;
  ram[25940]  = 1;
  ram[25941]  = 1;
  ram[25942]  = 1;
  ram[25943]  = 1;
  ram[25944]  = 1;
  ram[25945]  = 1;
  ram[25946]  = 1;
  ram[25947]  = 1;
  ram[25948]  = 1;
  ram[25949]  = 1;
  ram[25950]  = 1;
  ram[25951]  = 1;
  ram[25952]  = 1;
  ram[25953]  = 1;
  ram[25954]  = 1;
  ram[25955]  = 1;
  ram[25956]  = 1;
  ram[25957]  = 1;
  ram[25958]  = 1;
  ram[25959]  = 1;
  ram[25960]  = 1;
  ram[25961]  = 1;
  ram[25962]  = 1;
  ram[25963]  = 1;
  ram[25964]  = 1;
  ram[25965]  = 1;
  ram[25966]  = 1;
  ram[25967]  = 1;
  ram[25968]  = 1;
  ram[25969]  = 1;
  ram[25970]  = 1;
  ram[25971]  = 1;
  ram[25972]  = 1;
  ram[25973]  = 1;
  ram[25974]  = 1;
  ram[25975]  = 1;
  ram[25976]  = 1;
  ram[25977]  = 1;
  ram[25978]  = 1;
  ram[25979]  = 1;
  ram[25980]  = 1;
  ram[25981]  = 1;
  ram[25982]  = 1;
  ram[25983]  = 1;
  ram[25984]  = 1;
  ram[25985]  = 1;
  ram[25986]  = 1;
  ram[25987]  = 1;
  ram[25988]  = 1;
  ram[25989]  = 1;
  ram[25990]  = 1;
  ram[25991]  = 1;
  ram[25992]  = 1;
  ram[25993]  = 1;
  ram[25994]  = 1;
  ram[25995]  = 1;
  ram[25996]  = 1;
  ram[25997]  = 1;
  ram[25998]  = 1;
  ram[25999]  = 1;
  ram[26000]  = 1;
  ram[26001]  = 1;
  ram[26002]  = 1;
  ram[26003]  = 1;
  ram[26004]  = 1;
  ram[26005]  = 1;
  ram[26006]  = 1;
  ram[26007]  = 1;
  ram[26008]  = 1;
  ram[26009]  = 1;
  ram[26010]  = 1;
  ram[26011]  = 1;
  ram[26012]  = 1;
  ram[26013]  = 1;
  ram[26014]  = 1;
  ram[26015]  = 1;
  ram[26016]  = 1;
  ram[26017]  = 1;
  ram[26018]  = 1;
  ram[26019]  = 1;
  ram[26020]  = 1;
  ram[26021]  = 1;
  ram[26022]  = 1;
  ram[26023]  = 1;
  ram[26024]  = 1;
  ram[26025]  = 1;
  ram[26026]  = 1;
  ram[26027]  = 1;
  ram[26028]  = 1;
  ram[26029]  = 1;
  ram[26030]  = 1;
  ram[26031]  = 1;
  ram[26032]  = 1;
  ram[26033]  = 1;
  ram[26034]  = 1;
  ram[26035]  = 1;
  ram[26036]  = 1;
  ram[26037]  = 1;
  ram[26038]  = 1;
  ram[26039]  = 1;
  ram[26040]  = 1;
  ram[26041]  = 1;
  ram[26042]  = 1;
  ram[26043]  = 1;
  ram[26044]  = 1;
  ram[26045]  = 1;
  ram[26046]  = 1;
  ram[26047]  = 1;
  ram[26048]  = 1;
  ram[26049]  = 1;
  ram[26050]  = 1;
  ram[26051]  = 1;
  ram[26052]  = 1;
  ram[26053]  = 1;
  ram[26054]  = 1;
  ram[26055]  = 1;
  ram[26056]  = 1;
  ram[26057]  = 1;
  ram[26058]  = 1;
  ram[26059]  = 1;
  ram[26060]  = 1;
  ram[26061]  = 1;
  ram[26062]  = 1;
  ram[26063]  = 1;
  ram[26064]  = 1;
  ram[26065]  = 1;
  ram[26066]  = 1;
  ram[26067]  = 1;
  ram[26068]  = 1;
  ram[26069]  = 1;
  ram[26070]  = 1;
  ram[26071]  = 1;
  ram[26072]  = 1;
  ram[26073]  = 1;
  ram[26074]  = 1;
  ram[26075]  = 1;
  ram[26076]  = 1;
  ram[26077]  = 1;
  ram[26078]  = 1;
  ram[26079]  = 1;
  ram[26080]  = 1;
  ram[26081]  = 1;
  ram[26082]  = 1;
  ram[26083]  = 1;
  ram[26084]  = 1;
  ram[26085]  = 1;
  ram[26086]  = 1;
  ram[26087]  = 1;
  ram[26088]  = 1;
  ram[26089]  = 1;
  ram[26090]  = 1;
  ram[26091]  = 1;
  ram[26092]  = 1;
  ram[26093]  = 1;
  ram[26094]  = 1;
  ram[26095]  = 1;
  ram[26096]  = 1;
  ram[26097]  = 1;
  ram[26098]  = 1;
  ram[26099]  = 1;
  ram[26100]  = 1;
  ram[26101]  = 1;
  ram[26102]  = 1;
  ram[26103]  = 1;
  ram[26104]  = 1;
  ram[26105]  = 1;
  ram[26106]  = 1;
  ram[26107]  = 1;
  ram[26108]  = 1;
  ram[26109]  = 1;
  ram[26110]  = 1;
  ram[26111]  = 1;
  ram[26112]  = 1;
  ram[26113]  = 1;
  ram[26114]  = 1;
  ram[26115]  = 1;
  ram[26116]  = 1;
  ram[26117]  = 1;
  ram[26118]  = 1;
  ram[26119]  = 1;
  ram[26120]  = 1;
  ram[26121]  = 1;
  ram[26122]  = 1;
  ram[26123]  = 1;
  ram[26124]  = 1;
  ram[26125]  = 1;
  ram[26126]  = 1;
  ram[26127]  = 1;
  ram[26128]  = 1;
  ram[26129]  = 1;
  ram[26130]  = 1;
  ram[26131]  = 1;
  ram[26132]  = 1;
  ram[26133]  = 1;
  ram[26134]  = 1;
  ram[26135]  = 1;
  ram[26136]  = 1;
  ram[26137]  = 1;
  ram[26138]  = 1;
  ram[26139]  = 1;
  ram[26140]  = 1;
  ram[26141]  = 1;
  ram[26142]  = 1;
  ram[26143]  = 1;
  ram[26144]  = 1;
  ram[26145]  = 1;
  ram[26146]  = 1;
  ram[26147]  = 1;
  ram[26148]  = 1;
  ram[26149]  = 1;
  ram[26150]  = 1;
  ram[26151]  = 1;
  ram[26152]  = 1;
  ram[26153]  = 1;
  ram[26154]  = 1;
  ram[26155]  = 1;
  ram[26156]  = 1;
  ram[26157]  = 1;
  ram[26158]  = 1;
  ram[26159]  = 1;
  ram[26160]  = 1;
  ram[26161]  = 1;
  ram[26162]  = 1;
  ram[26163]  = 1;
  ram[26164]  = 1;
  ram[26165]  = 1;
  ram[26166]  = 1;
  ram[26167]  = 1;
  ram[26168]  = 1;
  ram[26169]  = 1;
  ram[26170]  = 1;
  ram[26171]  = 1;
  ram[26172]  = 1;
  ram[26173]  = 1;
  ram[26174]  = 1;
  ram[26175]  = 1;
  ram[26176]  = 1;
  ram[26177]  = 1;
  ram[26178]  = 1;
  ram[26179]  = 1;
  ram[26180]  = 1;
  ram[26181]  = 1;
  ram[26182]  = 1;
  ram[26183]  = 1;
  ram[26184]  = 1;
  ram[26185]  = 1;
  ram[26186]  = 1;
  ram[26187]  = 1;
  ram[26188]  = 1;
  ram[26189]  = 1;
  ram[26190]  = 1;
  ram[26191]  = 1;
  ram[26192]  = 1;
  ram[26193]  = 1;
  ram[26194]  = 1;
  ram[26195]  = 1;
  ram[26196]  = 1;
  ram[26197]  = 1;
  ram[26198]  = 1;
  ram[26199]  = 1;
  ram[26200]  = 1;
  ram[26201]  = 1;
  ram[26202]  = 1;
  ram[26203]  = 1;
  ram[26204]  = 1;
  ram[26205]  = 1;
  ram[26206]  = 1;
  ram[26207]  = 1;
  ram[26208]  = 1;
  ram[26209]  = 1;
  ram[26210]  = 1;
  ram[26211]  = 1;
  ram[26212]  = 1;
  ram[26213]  = 1;
  ram[26214]  = 1;
  ram[26215]  = 1;
  ram[26216]  = 1;
  ram[26217]  = 1;
  ram[26218]  = 1;
  ram[26219]  = 1;
  ram[26220]  = 1;
  ram[26221]  = 1;
  ram[26222]  = 1;
  ram[26223]  = 1;
  ram[26224]  = 1;
  ram[26225]  = 1;
  ram[26226]  = 1;
  ram[26227]  = 1;
  ram[26228]  = 1;
  ram[26229]  = 1;
  ram[26230]  = 1;
  ram[26231]  = 1;
  ram[26232]  = 1;
  ram[26233]  = 1;
  ram[26234]  = 1;
  ram[26235]  = 1;
  ram[26236]  = 1;
  ram[26237]  = 1;
  ram[26238]  = 1;
  ram[26239]  = 1;
  ram[26240]  = 1;
  ram[26241]  = 1;
  ram[26242]  = 1;
  ram[26243]  = 1;
  ram[26244]  = 1;
  ram[26245]  = 1;
  ram[26246]  = 1;
  ram[26247]  = 1;
  ram[26248]  = 1;
  ram[26249]  = 1;
  ram[26250]  = 1;
  ram[26251]  = 1;
  ram[26252]  = 1;
  ram[26253]  = 1;
  ram[26254]  = 1;
  ram[26255]  = 1;
  ram[26256]  = 1;
  ram[26257]  = 1;
  ram[26258]  = 1;
  ram[26259]  = 1;
  ram[26260]  = 1;
  ram[26261]  = 1;
  ram[26262]  = 1;
  ram[26263]  = 1;
  ram[26264]  = 1;
  ram[26265]  = 1;
  ram[26266]  = 1;
  ram[26267]  = 1;
  ram[26268]  = 1;
  ram[26269]  = 1;
  ram[26270]  = 1;
  ram[26271]  = 1;
  ram[26272]  = 1;
  ram[26273]  = 1;
  ram[26274]  = 1;
  ram[26275]  = 1;
  ram[26276]  = 1;
  ram[26277]  = 1;
  ram[26278]  = 1;
  ram[26279]  = 1;
  ram[26280]  = 1;
  ram[26281]  = 1;
  ram[26282]  = 1;
  ram[26283]  = 1;
  ram[26284]  = 1;
  ram[26285]  = 1;
  ram[26286]  = 1;
  ram[26287]  = 1;
  ram[26288]  = 1;
  ram[26289]  = 1;
  ram[26290]  = 1;
  ram[26291]  = 1;
  ram[26292]  = 1;
  ram[26293]  = 1;
  ram[26294]  = 1;
  ram[26295]  = 1;
  ram[26296]  = 1;
  ram[26297]  = 1;
  ram[26298]  = 1;
  ram[26299]  = 1;
  ram[26300]  = 1;
  ram[26301]  = 1;
  ram[26302]  = 1;
  ram[26303]  = 1;
  ram[26304]  = 1;
  ram[26305]  = 1;
  ram[26306]  = 1;
  ram[26307]  = 1;
  ram[26308]  = 1;
  ram[26309]  = 1;
  ram[26310]  = 1;
  ram[26311]  = 1;
  ram[26312]  = 1;
  ram[26313]  = 1;
  ram[26314]  = 1;
  ram[26315]  = 1;
  ram[26316]  = 1;
  ram[26317]  = 1;
  ram[26318]  = 1;
  ram[26319]  = 1;
  ram[26320]  = 1;
  ram[26321]  = 1;
  ram[26322]  = 1;
  ram[26323]  = 1;
  ram[26324]  = 1;
  ram[26325]  = 1;
  ram[26326]  = 1;
  ram[26327]  = 1;
  ram[26328]  = 1;
  ram[26329]  = 1;
  ram[26330]  = 1;
  ram[26331]  = 1;
  ram[26332]  = 1;
  ram[26333]  = 1;
  ram[26334]  = 1;
  ram[26335]  = 1;
  ram[26336]  = 1;
  ram[26337]  = 1;
  ram[26338]  = 1;
  ram[26339]  = 1;
  ram[26340]  = 1;
  ram[26341]  = 1;
  ram[26342]  = 1;
  ram[26343]  = 1;
  ram[26344]  = 1;
  ram[26345]  = 1;
  ram[26346]  = 1;
  ram[26347]  = 1;
  ram[26348]  = 1;
  ram[26349]  = 1;
  ram[26350]  = 1;
  ram[26351]  = 1;
  ram[26352]  = 1;
  ram[26353]  = 1;
  ram[26354]  = 1;
  ram[26355]  = 1;
  ram[26356]  = 1;
  ram[26357]  = 1;
  ram[26358]  = 1;
  ram[26359]  = 1;
  ram[26360]  = 1;
  ram[26361]  = 1;
  ram[26362]  = 1;
  ram[26363]  = 1;
  ram[26364]  = 1;
  ram[26365]  = 1;
  ram[26366]  = 1;
  ram[26367]  = 1;
  ram[26368]  = 1;
  ram[26369]  = 1;
  ram[26370]  = 1;
  ram[26371]  = 1;
  ram[26372]  = 1;
  ram[26373]  = 1;
  ram[26374]  = 1;
  ram[26375]  = 1;
  ram[26376]  = 1;
  ram[26377]  = 1;
  ram[26378]  = 1;
  ram[26379]  = 1;
  ram[26380]  = 1;
  ram[26381]  = 1;
  ram[26382]  = 1;
  ram[26383]  = 1;
  ram[26384]  = 1;
  ram[26385]  = 1;
  ram[26386]  = 1;
  ram[26387]  = 1;
  ram[26388]  = 1;
  ram[26389]  = 1;
  ram[26390]  = 1;
  ram[26391]  = 1;
  ram[26392]  = 1;
  ram[26393]  = 1;
  ram[26394]  = 1;
  ram[26395]  = 1;
  ram[26396]  = 1;
  ram[26397]  = 1;
  ram[26398]  = 1;
  ram[26399]  = 1;
  ram[26400]  = 1;
  ram[26401]  = 1;
  ram[26402]  = 1;
  ram[26403]  = 1;
  ram[26404]  = 1;
  ram[26405]  = 1;
  ram[26406]  = 1;
  ram[26407]  = 1;
  ram[26408]  = 1;
  ram[26409]  = 1;
  ram[26410]  = 1;
  ram[26411]  = 1;
  ram[26412]  = 1;
  ram[26413]  = 1;
  ram[26414]  = 1;
  ram[26415]  = 1;
  ram[26416]  = 1;
  ram[26417]  = 1;
  ram[26418]  = 1;
  ram[26419]  = 1;
  ram[26420]  = 1;
  ram[26421]  = 1;
  ram[26422]  = 1;
  ram[26423]  = 1;
  ram[26424]  = 1;
  ram[26425]  = 1;
  ram[26426]  = 1;
  ram[26427]  = 1;
  ram[26428]  = 1;
  ram[26429]  = 1;
  ram[26430]  = 1;
  ram[26431]  = 1;
  ram[26432]  = 1;
  ram[26433]  = 1;
  ram[26434]  = 1;
  ram[26435]  = 1;
  ram[26436]  = 1;
  ram[26437]  = 1;
  ram[26438]  = 1;
  ram[26439]  = 1;
  ram[26440]  = 1;
  ram[26441]  = 1;
  ram[26442]  = 1;
  ram[26443]  = 1;
  ram[26444]  = 1;
  ram[26445]  = 1;
  ram[26446]  = 1;
  ram[26447]  = 1;
  ram[26448]  = 1;
  ram[26449]  = 1;
  ram[26450]  = 1;
  ram[26451]  = 1;
  ram[26452]  = 1;
  ram[26453]  = 1;
  ram[26454]  = 1;
  ram[26455]  = 1;
  ram[26456]  = 1;
  ram[26457]  = 1;
  ram[26458]  = 1;
  ram[26459]  = 1;
  ram[26460]  = 1;
  ram[26461]  = 1;
  ram[26462]  = 1;
  ram[26463]  = 1;
  ram[26464]  = 1;
  ram[26465]  = 1;
  ram[26466]  = 1;
  ram[26467]  = 1;
  ram[26468]  = 1;
  ram[26469]  = 1;
  ram[26470]  = 1;
  ram[26471]  = 1;
  ram[26472]  = 1;
  ram[26473]  = 1;
  ram[26474]  = 1;
  ram[26475]  = 1;
  ram[26476]  = 1;
  ram[26477]  = 1;
  ram[26478]  = 1;
  ram[26479]  = 1;
  ram[26480]  = 1;
  ram[26481]  = 1;
  ram[26482]  = 1;
  ram[26483]  = 1;
  ram[26484]  = 1;
  ram[26485]  = 1;
  ram[26486]  = 1;
  ram[26487]  = 1;
  ram[26488]  = 1;
  ram[26489]  = 1;
  ram[26490]  = 1;
  ram[26491]  = 1;
  ram[26492]  = 1;
  ram[26493]  = 1;
  ram[26494]  = 1;
  ram[26495]  = 1;
  ram[26496]  = 1;
  ram[26497]  = 1;
  ram[26498]  = 1;
  ram[26499]  = 1;
  ram[26500]  = 1;
  ram[26501]  = 1;
  ram[26502]  = 1;
  ram[26503]  = 1;
  ram[26504]  = 1;
  ram[26505]  = 1;
  ram[26506]  = 1;
  ram[26507]  = 1;
  ram[26508]  = 1;
  ram[26509]  = 1;
  ram[26510]  = 1;
  ram[26511]  = 1;
  ram[26512]  = 1;
  ram[26513]  = 1;
  ram[26514]  = 1;
  ram[26515]  = 1;
  ram[26516]  = 1;
  ram[26517]  = 1;
  ram[26518]  = 1;
  ram[26519]  = 1;
  ram[26520]  = 1;
  ram[26521]  = 1;
  ram[26522]  = 1;
  ram[26523]  = 1;
  ram[26524]  = 1;
  ram[26525]  = 1;
  ram[26526]  = 1;
  ram[26527]  = 1;
  ram[26528]  = 1;
  ram[26529]  = 1;
  ram[26530]  = 1;
  ram[26531]  = 1;
  ram[26532]  = 1;
  ram[26533]  = 1;
  ram[26534]  = 1;
  ram[26535]  = 1;
  ram[26536]  = 1;
  ram[26537]  = 1;
  ram[26538]  = 1;
  ram[26539]  = 1;
  ram[26540]  = 1;
  ram[26541]  = 1;
  ram[26542]  = 1;
  ram[26543]  = 1;
  ram[26544]  = 1;
  ram[26545]  = 1;
  ram[26546]  = 1;
  ram[26547]  = 1;
  ram[26548]  = 1;
  ram[26549]  = 1;
  ram[26550]  = 1;
  ram[26551]  = 1;
  ram[26552]  = 1;
  ram[26553]  = 1;
  ram[26554]  = 1;
  ram[26555]  = 1;
  ram[26556]  = 1;
  ram[26557]  = 1;
  ram[26558]  = 1;
  ram[26559]  = 1;
  ram[26560]  = 1;
  ram[26561]  = 1;
  ram[26562]  = 1;
  ram[26563]  = 1;
  ram[26564]  = 1;
  ram[26565]  = 1;
  ram[26566]  = 1;
  ram[26567]  = 1;
  ram[26568]  = 1;
  ram[26569]  = 1;
  ram[26570]  = 1;
  ram[26571]  = 1;
  ram[26572]  = 1;
  ram[26573]  = 1;
  ram[26574]  = 1;
  ram[26575]  = 1;
  ram[26576]  = 1;
  ram[26577]  = 1;
  ram[26578]  = 1;
  ram[26579]  = 1;
  ram[26580]  = 1;
  ram[26581]  = 1;
  ram[26582]  = 1;
  ram[26583]  = 1;
  ram[26584]  = 1;
  ram[26585]  = 1;
  ram[26586]  = 1;
  ram[26587]  = 1;
  ram[26588]  = 1;
  ram[26589]  = 1;
  ram[26590]  = 1;
  ram[26591]  = 1;
  ram[26592]  = 1;
  ram[26593]  = 1;
  ram[26594]  = 1;
  ram[26595]  = 1;
  ram[26596]  = 1;
  ram[26597]  = 1;
  ram[26598]  = 1;
  ram[26599]  = 1;
  ram[26600]  = 1;
  ram[26601]  = 1;
  ram[26602]  = 1;
  ram[26603]  = 1;
  ram[26604]  = 1;
  ram[26605]  = 1;
  ram[26606]  = 1;
  ram[26607]  = 1;
  ram[26608]  = 1;
  ram[26609]  = 1;
  ram[26610]  = 1;
  ram[26611]  = 1;
  ram[26612]  = 1;
  ram[26613]  = 1;
  ram[26614]  = 1;
  ram[26615]  = 1;
  ram[26616]  = 1;
  ram[26617]  = 1;
  ram[26618]  = 1;
  ram[26619]  = 1;
  ram[26620]  = 1;
  ram[26621]  = 1;
  ram[26622]  = 1;
  ram[26623]  = 1;
  ram[26624]  = 1;
  ram[26625]  = 1;
  ram[26626]  = 1;
  ram[26627]  = 1;
  ram[26628]  = 1;
  ram[26629]  = 1;
  ram[26630]  = 1;
  ram[26631]  = 1;
  ram[26632]  = 1;
  ram[26633]  = 1;
  ram[26634]  = 1;
  ram[26635]  = 1;
  ram[26636]  = 1;
  ram[26637]  = 1;
  ram[26638]  = 1;
  ram[26639]  = 1;
  ram[26640]  = 1;
  ram[26641]  = 1;
  ram[26642]  = 1;
  ram[26643]  = 1;
  ram[26644]  = 1;
  ram[26645]  = 1;
  ram[26646]  = 1;
  ram[26647]  = 1;
  ram[26648]  = 1;
  ram[26649]  = 1;
  ram[26650]  = 1;
  ram[26651]  = 1;
  ram[26652]  = 1;
  ram[26653]  = 1;
  ram[26654]  = 1;
  ram[26655]  = 1;
  ram[26656]  = 1;
  ram[26657]  = 1;
  ram[26658]  = 1;
  ram[26659]  = 1;
  ram[26660]  = 1;
  ram[26661]  = 1;
  ram[26662]  = 1;
  ram[26663]  = 1;
  ram[26664]  = 1;
  ram[26665]  = 1;
  ram[26666]  = 1;
  ram[26667]  = 1;
  ram[26668]  = 1;
  ram[26669]  = 1;
  ram[26670]  = 1;
  ram[26671]  = 1;
  ram[26672]  = 1;
  ram[26673]  = 1;
  ram[26674]  = 1;
  ram[26675]  = 1;
  ram[26676]  = 1;
  ram[26677]  = 1;
  ram[26678]  = 1;
  ram[26679]  = 1;
  ram[26680]  = 1;
  ram[26681]  = 1;
  ram[26682]  = 1;
  ram[26683]  = 1;
  ram[26684]  = 1;
  ram[26685]  = 1;
  ram[26686]  = 1;
  ram[26687]  = 1;
  ram[26688]  = 1;
  ram[26689]  = 1;
  ram[26690]  = 1;
  ram[26691]  = 1;
  ram[26692]  = 1;
  ram[26693]  = 1;
  ram[26694]  = 1;
  ram[26695]  = 1;
  ram[26696]  = 1;
  ram[26697]  = 1;
  ram[26698]  = 1;
  ram[26699]  = 1;
  ram[26700]  = 1;
  ram[26701]  = 1;
  ram[26702]  = 1;
  ram[26703]  = 1;
  ram[26704]  = 1;
  ram[26705]  = 1;
  ram[26706]  = 1;
  ram[26707]  = 1;
  ram[26708]  = 1;
  ram[26709]  = 1;
  ram[26710]  = 1;
  ram[26711]  = 1;
  ram[26712]  = 1;
  ram[26713]  = 1;
  ram[26714]  = 1;
  ram[26715]  = 1;
  ram[26716]  = 1;
  ram[26717]  = 1;
  ram[26718]  = 1;
  ram[26719]  = 1;
  ram[26720]  = 1;
  ram[26721]  = 1;
  ram[26722]  = 1;
  ram[26723]  = 1;
  ram[26724]  = 1;
  ram[26725]  = 1;
  ram[26726]  = 1;
  ram[26727]  = 1;
  ram[26728]  = 1;
  ram[26729]  = 1;
  ram[26730]  = 1;
  ram[26731]  = 1;
  ram[26732]  = 1;
  ram[26733]  = 1;
  ram[26734]  = 1;
  ram[26735]  = 1;
  ram[26736]  = 1;
  ram[26737]  = 1;
  ram[26738]  = 1;
  ram[26739]  = 1;
  ram[26740]  = 1;
  ram[26741]  = 1;
  ram[26742]  = 1;
  ram[26743]  = 1;
  ram[26744]  = 1;
  ram[26745]  = 1;
  ram[26746]  = 1;
  ram[26747]  = 1;
  ram[26748]  = 1;
  ram[26749]  = 1;
  ram[26750]  = 1;
  ram[26751]  = 1;
  ram[26752]  = 1;
  ram[26753]  = 1;
  ram[26754]  = 1;
  ram[26755]  = 1;
  ram[26756]  = 1;
  ram[26757]  = 1;
  ram[26758]  = 1;
  ram[26759]  = 1;
  ram[26760]  = 1;
  ram[26761]  = 1;
  ram[26762]  = 1;
  ram[26763]  = 1;
  ram[26764]  = 1;
  ram[26765]  = 1;
  ram[26766]  = 1;
  ram[26767]  = 1;
  ram[26768]  = 1;
  ram[26769]  = 1;
  ram[26770]  = 1;
  ram[26771]  = 1;
  ram[26772]  = 1;
  ram[26773]  = 1;
  ram[26774]  = 1;
  ram[26775]  = 1;
  ram[26776]  = 1;
  ram[26777]  = 1;
  ram[26778]  = 1;
  ram[26779]  = 1;
  ram[26780]  = 1;
  ram[26781]  = 1;
  ram[26782]  = 1;
  ram[26783]  = 1;
  ram[26784]  = 1;
  ram[26785]  = 1;
  ram[26786]  = 1;
  ram[26787]  = 1;
  ram[26788]  = 1;
  ram[26789]  = 1;
  ram[26790]  = 1;
  ram[26791]  = 1;
  ram[26792]  = 1;
  ram[26793]  = 1;
  ram[26794]  = 1;
  ram[26795]  = 1;
  ram[26796]  = 1;
  ram[26797]  = 1;
  ram[26798]  = 1;
  ram[26799]  = 1;
  ram[26800]  = 1;
  ram[26801]  = 1;
  ram[26802]  = 1;
  ram[26803]  = 1;
  ram[26804]  = 1;
  ram[26805]  = 1;
  ram[26806]  = 1;
  ram[26807]  = 1;
  ram[26808]  = 1;
  ram[26809]  = 1;
  ram[26810]  = 1;
  ram[26811]  = 1;
  ram[26812]  = 1;
  ram[26813]  = 1;
  ram[26814]  = 1;
  ram[26815]  = 1;
  ram[26816]  = 1;
  ram[26817]  = 1;
  ram[26818]  = 1;
  ram[26819]  = 1;
  ram[26820]  = 1;
  ram[26821]  = 1;
  ram[26822]  = 1;
  ram[26823]  = 1;
  ram[26824]  = 1;
  ram[26825]  = 1;
  ram[26826]  = 1;
  ram[26827]  = 1;
  ram[26828]  = 1;
  ram[26829]  = 1;
  ram[26830]  = 1;
  ram[26831]  = 1;
  ram[26832]  = 1;
  ram[26833]  = 1;
  ram[26834]  = 1;
  ram[26835]  = 1;
  ram[26836]  = 1;
  ram[26837]  = 1;
  ram[26838]  = 1;
  ram[26839]  = 1;
  ram[26840]  = 1;
  ram[26841]  = 1;
  ram[26842]  = 1;
  ram[26843]  = 1;
  ram[26844]  = 1;
  ram[26845]  = 1;
  ram[26846]  = 1;
  ram[26847]  = 1;
  ram[26848]  = 1;
  ram[26849]  = 1;
  ram[26850]  = 1;
  ram[26851]  = 1;
  ram[26852]  = 1;
  ram[26853]  = 1;
  ram[26854]  = 1;
  ram[26855]  = 1;
  ram[26856]  = 1;
  ram[26857]  = 1;
  ram[26858]  = 1;
  ram[26859]  = 1;
  ram[26860]  = 1;
  ram[26861]  = 1;
  ram[26862]  = 1;
  ram[26863]  = 1;
  ram[26864]  = 1;
  ram[26865]  = 1;
  ram[26866]  = 1;
  ram[26867]  = 1;
  ram[26868]  = 1;
  ram[26869]  = 1;
  ram[26870]  = 1;
  ram[26871]  = 1;
  ram[26872]  = 1;
  ram[26873]  = 1;
  ram[26874]  = 1;
  ram[26875]  = 1;
  ram[26876]  = 1;
  ram[26877]  = 1;
  ram[26878]  = 1;
  ram[26879]  = 1;
  ram[26880]  = 1;
  ram[26881]  = 1;
  ram[26882]  = 1;
  ram[26883]  = 1;
  ram[26884]  = 1;
  ram[26885]  = 1;
  ram[26886]  = 1;
  ram[26887]  = 1;
  ram[26888]  = 1;
  ram[26889]  = 1;
  ram[26890]  = 1;
  ram[26891]  = 1;
  ram[26892]  = 1;
  ram[26893]  = 1;
  ram[26894]  = 1;
  ram[26895]  = 1;
  ram[26896]  = 1;
  ram[26897]  = 1;
  ram[26898]  = 1;
  ram[26899]  = 1;
  ram[26900]  = 1;
  ram[26901]  = 1;
  ram[26902]  = 1;
  ram[26903]  = 1;
  ram[26904]  = 1;
  ram[26905]  = 1;
  ram[26906]  = 1;
  ram[26907]  = 1;
  ram[26908]  = 1;
  ram[26909]  = 1;
  ram[26910]  = 1;
  ram[26911]  = 1;
  ram[26912]  = 1;
  ram[26913]  = 1;
  ram[26914]  = 1;
  ram[26915]  = 1;
  ram[26916]  = 1;
  ram[26917]  = 1;
  ram[26918]  = 1;
  ram[26919]  = 1;
  ram[26920]  = 1;
  ram[26921]  = 1;
  ram[26922]  = 1;
  ram[26923]  = 1;
  ram[26924]  = 1;
  ram[26925]  = 1;
  ram[26926]  = 1;
  ram[26927]  = 1;
  ram[26928]  = 1;
  ram[26929]  = 1;
  ram[26930]  = 1;
  ram[26931]  = 1;
  ram[26932]  = 1;
  ram[26933]  = 1;
  ram[26934]  = 1;
  ram[26935]  = 1;
  ram[26936]  = 1;
  ram[26937]  = 1;
  ram[26938]  = 1;
  ram[26939]  = 1;
  ram[26940]  = 1;
  ram[26941]  = 1;
  ram[26942]  = 1;
  ram[26943]  = 1;
  ram[26944]  = 1;
  ram[26945]  = 1;
  ram[26946]  = 1;
  ram[26947]  = 1;
  ram[26948]  = 1;
  ram[26949]  = 1;
  ram[26950]  = 1;
  ram[26951]  = 1;
  ram[26952]  = 1;
  ram[26953]  = 1;
  ram[26954]  = 1;
  ram[26955]  = 1;
  ram[26956]  = 1;
  ram[26957]  = 1;
  ram[26958]  = 1;
  ram[26959]  = 1;
  ram[26960]  = 1;
  ram[26961]  = 1;
  ram[26962]  = 1;
  ram[26963]  = 1;
  ram[26964]  = 1;
  ram[26965]  = 1;
  ram[26966]  = 1;
  ram[26967]  = 1;
  ram[26968]  = 1;
  ram[26969]  = 1;
  ram[26970]  = 1;
  ram[26971]  = 1;
  ram[26972]  = 1;
  ram[26973]  = 1;
  ram[26974]  = 1;
  ram[26975]  = 1;
  ram[26976]  = 1;
  ram[26977]  = 1;
  ram[26978]  = 1;
  ram[26979]  = 1;
  ram[26980]  = 1;
  ram[26981]  = 1;
  ram[26982]  = 1;
  ram[26983]  = 1;
  ram[26984]  = 1;
  ram[26985]  = 1;
  ram[26986]  = 1;
  ram[26987]  = 1;
  ram[26988]  = 1;
  ram[26989]  = 1;
  ram[26990]  = 1;
  ram[26991]  = 1;
  ram[26992]  = 1;
  ram[26993]  = 1;
  ram[26994]  = 1;
  ram[26995]  = 1;
  ram[26996]  = 1;
  ram[26997]  = 1;
  ram[26998]  = 1;
  ram[26999]  = 1;
  ram[27000]  = 1;
  ram[27001]  = 1;
  ram[27002]  = 1;
  ram[27003]  = 1;
  ram[27004]  = 1;
  ram[27005]  = 1;
  ram[27006]  = 1;
  ram[27007]  = 1;
  ram[27008]  = 1;
  ram[27009]  = 1;
  ram[27010]  = 1;
  ram[27011]  = 1;
  ram[27012]  = 1;
  ram[27013]  = 1;
  ram[27014]  = 1;
  ram[27015]  = 1;
  ram[27016]  = 1;
  ram[27017]  = 1;
  ram[27018]  = 1;
  ram[27019]  = 1;
  ram[27020]  = 1;
  ram[27021]  = 1;
  ram[27022]  = 1;
  ram[27023]  = 1;
  ram[27024]  = 1;
  ram[27025]  = 1;
  ram[27026]  = 1;
  ram[27027]  = 1;
  ram[27028]  = 1;
  ram[27029]  = 1;
  ram[27030]  = 1;
  ram[27031]  = 1;
  ram[27032]  = 1;
  ram[27033]  = 1;
  ram[27034]  = 1;
  ram[27035]  = 1;
  ram[27036]  = 1;
  ram[27037]  = 1;
  ram[27038]  = 1;
  ram[27039]  = 1;
  ram[27040]  = 1;
  ram[27041]  = 1;
  ram[27042]  = 1;
  ram[27043]  = 1;
  ram[27044]  = 1;
  ram[27045]  = 1;
  ram[27046]  = 1;
  ram[27047]  = 1;
  ram[27048]  = 1;
  ram[27049]  = 1;
  ram[27050]  = 1;
  ram[27051]  = 1;
  ram[27052]  = 1;
  ram[27053]  = 1;
  ram[27054]  = 1;
  ram[27055]  = 1;
  ram[27056]  = 1;
  ram[27057]  = 1;
  ram[27058]  = 1;
  ram[27059]  = 1;
  ram[27060]  = 1;
  ram[27061]  = 1;
  ram[27062]  = 1;
  ram[27063]  = 1;
  ram[27064]  = 1;
  ram[27065]  = 1;
  ram[27066]  = 1;
  ram[27067]  = 1;
  ram[27068]  = 1;
  ram[27069]  = 1;
  ram[27070]  = 1;
  ram[27071]  = 1;
  ram[27072]  = 1;
  ram[27073]  = 1;
  ram[27074]  = 1;
  ram[27075]  = 1;
  ram[27076]  = 1;
  ram[27077]  = 1;
  ram[27078]  = 1;
  ram[27079]  = 1;
  ram[27080]  = 1;
  ram[27081]  = 1;
  ram[27082]  = 1;
  ram[27083]  = 1;
  ram[27084]  = 1;
  ram[27085]  = 1;
  ram[27086]  = 1;
  ram[27087]  = 1;
  ram[27088]  = 1;
  ram[27089]  = 1;
  ram[27090]  = 1;
  ram[27091]  = 1;
  ram[27092]  = 1;
  ram[27093]  = 1;
  ram[27094]  = 1;
  ram[27095]  = 1;
  ram[27096]  = 1;
  ram[27097]  = 1;
  ram[27098]  = 1;
  ram[27099]  = 1;
  ram[27100]  = 1;
  ram[27101]  = 1;
  ram[27102]  = 1;
  ram[27103]  = 1;
  ram[27104]  = 1;
  ram[27105]  = 1;
  ram[27106]  = 1;
  ram[27107]  = 1;
  ram[27108]  = 1;
  ram[27109]  = 1;
  ram[27110]  = 1;
  ram[27111]  = 1;
  ram[27112]  = 1;
  ram[27113]  = 1;
  ram[27114]  = 1;
  ram[27115]  = 1;
  ram[27116]  = 1;
  ram[27117]  = 1;
  ram[27118]  = 1;
  ram[27119]  = 1;
  ram[27120]  = 1;
  ram[27121]  = 1;
  ram[27122]  = 1;
  ram[27123]  = 1;
  ram[27124]  = 1;
  ram[27125]  = 1;
  ram[27126]  = 1;
  ram[27127]  = 1;
  ram[27128]  = 1;
  ram[27129]  = 1;
  ram[27130]  = 1;
  ram[27131]  = 1;
  ram[27132]  = 1;
  ram[27133]  = 1;
  ram[27134]  = 1;
  ram[27135]  = 1;
  ram[27136]  = 1;
  ram[27137]  = 1;
  ram[27138]  = 1;
  ram[27139]  = 1;
  ram[27140]  = 1;
  ram[27141]  = 1;
  ram[27142]  = 1;
  ram[27143]  = 1;
  ram[27144]  = 1;
  ram[27145]  = 1;
  ram[27146]  = 1;
  ram[27147]  = 1;
  ram[27148]  = 1;
  ram[27149]  = 1;
  ram[27150]  = 1;
  ram[27151]  = 1;
  ram[27152]  = 1;
  ram[27153]  = 1;
  ram[27154]  = 1;
  ram[27155]  = 1;
  ram[27156]  = 1;
  ram[27157]  = 1;
  ram[27158]  = 1;
  ram[27159]  = 1;
  ram[27160]  = 1;
  ram[27161]  = 1;
  ram[27162]  = 1;
  ram[27163]  = 1;
  ram[27164]  = 1;
  ram[27165]  = 1;
  ram[27166]  = 1;
  ram[27167]  = 1;
  ram[27168]  = 1;
  ram[27169]  = 1;
  ram[27170]  = 1;
  ram[27171]  = 1;
  ram[27172]  = 1;
  ram[27173]  = 1;
  ram[27174]  = 1;
  ram[27175]  = 1;
  ram[27176]  = 1;
  ram[27177]  = 1;
  ram[27178]  = 1;
  ram[27179]  = 1;
  ram[27180]  = 1;
  ram[27181]  = 1;
  ram[27182]  = 1;
  ram[27183]  = 1;
  ram[27184]  = 1;
  ram[27185]  = 1;
  ram[27186]  = 1;
  ram[27187]  = 1;
  ram[27188]  = 1;
  ram[27189]  = 1;
  ram[27190]  = 1;
  ram[27191]  = 1;
  ram[27192]  = 1;
  ram[27193]  = 1;
  ram[27194]  = 1;
  ram[27195]  = 1;
  ram[27196]  = 1;
  ram[27197]  = 1;
  ram[27198]  = 1;
  ram[27199]  = 1;
  ram[27200]  = 1;
  ram[27201]  = 1;
  ram[27202]  = 1;
  ram[27203]  = 1;
  ram[27204]  = 1;
  ram[27205]  = 1;
  ram[27206]  = 1;
  ram[27207]  = 1;
  ram[27208]  = 1;
  ram[27209]  = 1;
  ram[27210]  = 1;
  ram[27211]  = 1;
  ram[27212]  = 1;
  ram[27213]  = 1;
  ram[27214]  = 1;
  ram[27215]  = 1;
  ram[27216]  = 1;
  ram[27217]  = 1;
  ram[27218]  = 1;
  ram[27219]  = 1;
  ram[27220]  = 1;
  ram[27221]  = 1;
  ram[27222]  = 1;
  ram[27223]  = 1;
  ram[27224]  = 1;
  ram[27225]  = 1;
  ram[27226]  = 1;
  ram[27227]  = 1;
  ram[27228]  = 1;
  ram[27229]  = 1;
  ram[27230]  = 1;
  ram[27231]  = 1;
  ram[27232]  = 1;
  ram[27233]  = 1;
  ram[27234]  = 1;
  ram[27235]  = 1;
  ram[27236]  = 1;
  ram[27237]  = 1;
  ram[27238]  = 1;
  ram[27239]  = 1;
  ram[27240]  = 1;
  ram[27241]  = 1;
  ram[27242]  = 1;
  ram[27243]  = 1;
  ram[27244]  = 1;
  ram[27245]  = 1;
  ram[27246]  = 1;
  ram[27247]  = 1;
  ram[27248]  = 1;
  ram[27249]  = 1;
  ram[27250]  = 1;
  ram[27251]  = 1;
  ram[27252]  = 1;
  ram[27253]  = 1;
  ram[27254]  = 1;
  ram[27255]  = 1;
  ram[27256]  = 1;
  ram[27257]  = 1;
  ram[27258]  = 1;
  ram[27259]  = 1;
  ram[27260]  = 1;
  ram[27261]  = 1;
  ram[27262]  = 1;
  ram[27263]  = 1;
  ram[27264]  = 1;
  ram[27265]  = 1;
  ram[27266]  = 1;
  ram[27267]  = 1;
  ram[27268]  = 1;
  ram[27269]  = 1;
  ram[27270]  = 1;
  ram[27271]  = 1;
  ram[27272]  = 1;
  ram[27273]  = 1;
  ram[27274]  = 1;
  ram[27275]  = 1;
  ram[27276]  = 1;
  ram[27277]  = 1;
  ram[27278]  = 1;
  ram[27279]  = 1;
  ram[27280]  = 1;
  ram[27281]  = 1;
  ram[27282]  = 1;
  ram[27283]  = 1;
  ram[27284]  = 1;
  ram[27285]  = 1;
  ram[27286]  = 1;
  ram[27287]  = 1;
  ram[27288]  = 1;
  ram[27289]  = 1;
  ram[27290]  = 1;
  ram[27291]  = 1;
  ram[27292]  = 1;
  ram[27293]  = 1;
  ram[27294]  = 1;
  ram[27295]  = 1;
  ram[27296]  = 1;
  ram[27297]  = 1;
  ram[27298]  = 1;
  ram[27299]  = 1;
  ram[27300]  = 1;
  ram[27301]  = 1;
  ram[27302]  = 1;
  ram[27303]  = 1;
  ram[27304]  = 1;
  ram[27305]  = 1;
  ram[27306]  = 1;
  ram[27307]  = 1;
  ram[27308]  = 1;
  ram[27309]  = 1;
  ram[27310]  = 1;
  ram[27311]  = 1;
  ram[27312]  = 1;
  ram[27313]  = 1;
  ram[27314]  = 1;
  ram[27315]  = 1;
  ram[27316]  = 1;
  ram[27317]  = 1;
  ram[27318]  = 1;
  ram[27319]  = 1;
  ram[27320]  = 1;
  ram[27321]  = 1;
  ram[27322]  = 1;
  ram[27323]  = 1;
  ram[27324]  = 1;
  ram[27325]  = 1;
  ram[27326]  = 1;
  ram[27327]  = 1;
  ram[27328]  = 1;
  ram[27329]  = 1;
  ram[27330]  = 1;
  ram[27331]  = 1;
  ram[27332]  = 1;
  ram[27333]  = 1;
  ram[27334]  = 1;
  ram[27335]  = 1;
  ram[27336]  = 1;
  ram[27337]  = 1;
  ram[27338]  = 1;
  ram[27339]  = 1;
  ram[27340]  = 1;
  ram[27341]  = 1;
  ram[27342]  = 1;
  ram[27343]  = 1;
  ram[27344]  = 1;
  ram[27345]  = 1;
  ram[27346]  = 1;
  ram[27347]  = 1;
  ram[27348]  = 1;
  ram[27349]  = 1;
  ram[27350]  = 1;
  ram[27351]  = 1;
  ram[27352]  = 1;
  ram[27353]  = 1;
  ram[27354]  = 1;
  ram[27355]  = 1;
  ram[27356]  = 1;
  ram[27357]  = 1;
  ram[27358]  = 1;
  ram[27359]  = 1;
  ram[27360]  = 1;
  ram[27361]  = 1;
  ram[27362]  = 1;
  ram[27363]  = 1;
  ram[27364]  = 1;
  ram[27365]  = 1;
  ram[27366]  = 1;
  ram[27367]  = 1;
  ram[27368]  = 1;
  ram[27369]  = 1;
  ram[27370]  = 1;
  ram[27371]  = 1;
  ram[27372]  = 1;
  ram[27373]  = 1;
  ram[27374]  = 1;
  ram[27375]  = 1;
  ram[27376]  = 1;
  ram[27377]  = 1;
  ram[27378]  = 1;
  ram[27379]  = 1;
  ram[27380]  = 1;
  ram[27381]  = 1;
  ram[27382]  = 1;
  ram[27383]  = 1;
  ram[27384]  = 1;
  ram[27385]  = 1;
  ram[27386]  = 1;
  ram[27387]  = 1;
  ram[27388]  = 1;
  ram[27389]  = 1;
  ram[27390]  = 1;
  ram[27391]  = 1;
  ram[27392]  = 1;
  ram[27393]  = 1;
  ram[27394]  = 1;
  ram[27395]  = 1;
  ram[27396]  = 1;
  ram[27397]  = 1;
  ram[27398]  = 1;
  ram[27399]  = 1;
  ram[27400]  = 1;
  ram[27401]  = 1;
  ram[27402]  = 1;
  ram[27403]  = 1;
  ram[27404]  = 1;
  ram[27405]  = 1;
  ram[27406]  = 1;
  ram[27407]  = 1;
  ram[27408]  = 1;
  ram[27409]  = 1;
  ram[27410]  = 1;
  ram[27411]  = 1;
  ram[27412]  = 1;
  ram[27413]  = 1;
  ram[27414]  = 1;
  ram[27415]  = 1;
  ram[27416]  = 1;
  ram[27417]  = 1;
  ram[27418]  = 1;
  ram[27419]  = 1;
  ram[27420]  = 1;
  ram[27421]  = 1;
  ram[27422]  = 1;
  ram[27423]  = 1;
  ram[27424]  = 1;
  ram[27425]  = 1;
  ram[27426]  = 1;
  ram[27427]  = 1;
  ram[27428]  = 1;
  ram[27429]  = 1;
  ram[27430]  = 1;
  ram[27431]  = 1;
  ram[27432]  = 1;
  ram[27433]  = 1;
  ram[27434]  = 1;
  ram[27435]  = 1;
  ram[27436]  = 1;
  ram[27437]  = 1;
  ram[27438]  = 1;
  ram[27439]  = 1;
  ram[27440]  = 1;
  ram[27441]  = 1;
  ram[27442]  = 1;
  ram[27443]  = 1;
  ram[27444]  = 1;
  ram[27445]  = 1;
  ram[27446]  = 1;
  ram[27447]  = 1;
  ram[27448]  = 1;
  ram[27449]  = 1;
  ram[27450]  = 1;
  ram[27451]  = 1;
  ram[27452]  = 1;
  ram[27453]  = 1;
  ram[27454]  = 1;
  ram[27455]  = 1;
  ram[27456]  = 1;
  ram[27457]  = 1;
  ram[27458]  = 1;
  ram[27459]  = 1;
  ram[27460]  = 1;
  ram[27461]  = 1;
  ram[27462]  = 1;
  ram[27463]  = 1;
  ram[27464]  = 1;
  ram[27465]  = 1;
  ram[27466]  = 1;
  ram[27467]  = 1;
  ram[27468]  = 1;
  ram[27469]  = 1;
  ram[27470]  = 1;
  ram[27471]  = 1;
  ram[27472]  = 1;
  ram[27473]  = 1;
  ram[27474]  = 1;
  ram[27475]  = 1;
  ram[27476]  = 1;
  ram[27477]  = 1;
  ram[27478]  = 1;
  ram[27479]  = 1;
  ram[27480]  = 1;
  ram[27481]  = 1;
  ram[27482]  = 1;
  ram[27483]  = 1;
  ram[27484]  = 1;
  ram[27485]  = 1;
  ram[27486]  = 1;
  ram[27487]  = 1;
  ram[27488]  = 1;
  ram[27489]  = 1;
  ram[27490]  = 1;
  ram[27491]  = 1;
  ram[27492]  = 1;
  ram[27493]  = 1;
  ram[27494]  = 1;
  ram[27495]  = 1;
  ram[27496]  = 1;
  ram[27497]  = 1;
  ram[27498]  = 1;
  ram[27499]  = 1;
  ram[27500]  = 1;
  ram[27501]  = 1;
  ram[27502]  = 1;
  ram[27503]  = 1;
  ram[27504]  = 1;
  ram[27505]  = 1;
  ram[27506]  = 1;
  ram[27507]  = 1;
  ram[27508]  = 1;
  ram[27509]  = 1;
  ram[27510]  = 1;
  ram[27511]  = 1;
  ram[27512]  = 1;
  ram[27513]  = 1;
  ram[27514]  = 1;
  ram[27515]  = 1;
  ram[27516]  = 1;
  ram[27517]  = 1;
  ram[27518]  = 1;
  ram[27519]  = 1;
  ram[27520]  = 1;
  ram[27521]  = 1;
  ram[27522]  = 1;
  ram[27523]  = 1;
  ram[27524]  = 1;
  ram[27525]  = 1;
  ram[27526]  = 1;
  ram[27527]  = 1;
  ram[27528]  = 1;
  ram[27529]  = 1;
  ram[27530]  = 1;
  ram[27531]  = 1;
  ram[27532]  = 1;
  ram[27533]  = 1;
  ram[27534]  = 1;
  ram[27535]  = 1;
  ram[27536]  = 1;
  ram[27537]  = 1;
  ram[27538]  = 1;
  ram[27539]  = 1;
  ram[27540]  = 1;
  ram[27541]  = 1;
  ram[27542]  = 1;
  ram[27543]  = 1;
  ram[27544]  = 1;
  ram[27545]  = 1;
  ram[27546]  = 1;
  ram[27547]  = 1;
  ram[27548]  = 1;
  ram[27549]  = 1;
  ram[27550]  = 1;
  ram[27551]  = 1;
  ram[27552]  = 1;
  ram[27553]  = 1;
  ram[27554]  = 1;
  ram[27555]  = 1;
  ram[27556]  = 1;
  ram[27557]  = 1;
  ram[27558]  = 1;
  ram[27559]  = 1;
  ram[27560]  = 1;
  ram[27561]  = 1;
  ram[27562]  = 1;
  ram[27563]  = 1;
  ram[27564]  = 1;
  ram[27565]  = 1;
  ram[27566]  = 1;
  ram[27567]  = 1;
  ram[27568]  = 1;
  ram[27569]  = 1;
  ram[27570]  = 1;
  ram[27571]  = 1;
  ram[27572]  = 1;
  ram[27573]  = 1;
  ram[27574]  = 1;
  ram[27575]  = 1;
  ram[27576]  = 1;
  ram[27577]  = 1;
  ram[27578]  = 1;
  ram[27579]  = 1;
  ram[27580]  = 1;
  ram[27581]  = 1;
  ram[27582]  = 1;
  ram[27583]  = 1;
  ram[27584]  = 1;
  ram[27585]  = 1;
  ram[27586]  = 1;
  ram[27587]  = 1;
  ram[27588]  = 1;
  ram[27589]  = 1;
  ram[27590]  = 1;
  ram[27591]  = 1;
  ram[27592]  = 1;
  ram[27593]  = 1;
  ram[27594]  = 1;
  ram[27595]  = 1;
  ram[27596]  = 1;
  ram[27597]  = 1;
  ram[27598]  = 1;
  ram[27599]  = 1;
  ram[27600]  = 1;
  ram[27601]  = 1;
  ram[27602]  = 1;
  ram[27603]  = 1;
  ram[27604]  = 1;
  ram[27605]  = 1;
  ram[27606]  = 1;
  ram[27607]  = 1;
  ram[27608]  = 1;
  ram[27609]  = 1;
  ram[27610]  = 1;
  ram[27611]  = 1;
  ram[27612]  = 1;
  ram[27613]  = 1;
  ram[27614]  = 1;
  ram[27615]  = 1;
  ram[27616]  = 1;
  ram[27617]  = 1;
  ram[27618]  = 1;
  ram[27619]  = 1;
  ram[27620]  = 1;
  ram[27621]  = 1;
  ram[27622]  = 1;
  ram[27623]  = 1;
  ram[27624]  = 1;
  ram[27625]  = 1;
  ram[27626]  = 1;
  ram[27627]  = 1;
  ram[27628]  = 1;
  ram[27629]  = 1;
  ram[27630]  = 1;
  ram[27631]  = 1;
  ram[27632]  = 1;
  ram[27633]  = 1;
  ram[27634]  = 1;
  ram[27635]  = 1;
  ram[27636]  = 1;
  ram[27637]  = 1;
  ram[27638]  = 1;
  ram[27639]  = 1;
  ram[27640]  = 1;
  ram[27641]  = 1;
  ram[27642]  = 1;
  ram[27643]  = 1;
  ram[27644]  = 1;
  ram[27645]  = 1;
  ram[27646]  = 1;
  ram[27647]  = 1;
  ram[27648]  = 1;
  ram[27649]  = 1;
  ram[27650]  = 1;
  ram[27651]  = 1;
  ram[27652]  = 1;
  ram[27653]  = 1;
  ram[27654]  = 1;
  ram[27655]  = 1;
  ram[27656]  = 1;
  ram[27657]  = 1;
  ram[27658]  = 1;
  ram[27659]  = 1;
  ram[27660]  = 1;
  ram[27661]  = 1;
  ram[27662]  = 1;
  ram[27663]  = 1;
  ram[27664]  = 1;
  ram[27665]  = 1;
  ram[27666]  = 1;
  ram[27667]  = 1;
  ram[27668]  = 1;
  ram[27669]  = 1;
  ram[27670]  = 1;
  ram[27671]  = 1;
  ram[27672]  = 1;
  ram[27673]  = 1;
  ram[27674]  = 1;
  ram[27675]  = 1;
  ram[27676]  = 1;
  ram[27677]  = 1;
  ram[27678]  = 1;
  ram[27679]  = 1;
  ram[27680]  = 1;
  ram[27681]  = 1;
  ram[27682]  = 1;
  ram[27683]  = 1;
  ram[27684]  = 1;
  ram[27685]  = 1;
  ram[27686]  = 1;
  ram[27687]  = 1;
  ram[27688]  = 1;
  ram[27689]  = 1;
  ram[27690]  = 1;
  ram[27691]  = 1;
  ram[27692]  = 1;
  ram[27693]  = 1;
  ram[27694]  = 1;
  ram[27695]  = 1;
  ram[27696]  = 1;
  ram[27697]  = 1;
  ram[27698]  = 1;
  ram[27699]  = 1;
  ram[27700]  = 1;
  ram[27701]  = 1;
  ram[27702]  = 1;
  ram[27703]  = 1;
  ram[27704]  = 1;
  ram[27705]  = 1;
  ram[27706]  = 1;
  ram[27707]  = 1;
  ram[27708]  = 1;
  ram[27709]  = 1;
  ram[27710]  = 1;
  ram[27711]  = 1;
  ram[27712]  = 1;
  ram[27713]  = 1;
  ram[27714]  = 1;
  ram[27715]  = 1;
  ram[27716]  = 1;
  ram[27717]  = 1;
  ram[27718]  = 1;
  ram[27719]  = 1;
  ram[27720]  = 1;
  ram[27721]  = 1;
  ram[27722]  = 1;
  ram[27723]  = 1;
  ram[27724]  = 1;
  ram[27725]  = 1;
  ram[27726]  = 1;
  ram[27727]  = 1;
  ram[27728]  = 1;
  ram[27729]  = 1;
  ram[27730]  = 1;
  ram[27731]  = 1;
  ram[27732]  = 1;
  ram[27733]  = 1;
  ram[27734]  = 1;
  ram[27735]  = 1;
  ram[27736]  = 1;
  ram[27737]  = 1;
  ram[27738]  = 1;
  ram[27739]  = 1;
  ram[27740]  = 1;
  ram[27741]  = 1;
  ram[27742]  = 1;
  ram[27743]  = 1;
  ram[27744]  = 1;
  ram[27745]  = 1;
  ram[27746]  = 1;
  ram[27747]  = 1;
  ram[27748]  = 1;
  ram[27749]  = 1;
  ram[27750]  = 1;
  ram[27751]  = 1;
  ram[27752]  = 1;
  ram[27753]  = 1;
  ram[27754]  = 1;
  ram[27755]  = 1;
  ram[27756]  = 1;
  ram[27757]  = 1;
  ram[27758]  = 1;
  ram[27759]  = 1;
  ram[27760]  = 1;
  ram[27761]  = 1;
  ram[27762]  = 1;
  ram[27763]  = 1;
  ram[27764]  = 1;
  ram[27765]  = 1;
  ram[27766]  = 1;
  ram[27767]  = 1;
  ram[27768]  = 1;
  ram[27769]  = 1;
  ram[27770]  = 1;
  ram[27771]  = 1;
  ram[27772]  = 1;
  ram[27773]  = 1;
  ram[27774]  = 1;
  ram[27775]  = 1;
  ram[27776]  = 1;
  ram[27777]  = 1;
  ram[27778]  = 1;
  ram[27779]  = 1;
  ram[27780]  = 1;
  ram[27781]  = 1;
  ram[27782]  = 1;
  ram[27783]  = 1;
  ram[27784]  = 1;
  ram[27785]  = 1;
  ram[27786]  = 1;
  ram[27787]  = 1;
  ram[27788]  = 1;
  ram[27789]  = 1;
  ram[27790]  = 1;
  ram[27791]  = 1;
  ram[27792]  = 1;
  ram[27793]  = 1;
  ram[27794]  = 1;
  ram[27795]  = 1;
  ram[27796]  = 1;
  ram[27797]  = 1;
  ram[27798]  = 1;
  ram[27799]  = 1;
  ram[27800]  = 1;
  ram[27801]  = 1;
  ram[27802]  = 1;
  ram[27803]  = 1;
  ram[27804]  = 1;
  ram[27805]  = 1;
  ram[27806]  = 1;
  ram[27807]  = 1;
  ram[27808]  = 1;
  ram[27809]  = 1;
  ram[27810]  = 1;
  ram[27811]  = 1;
  ram[27812]  = 1;
  ram[27813]  = 1;
  ram[27814]  = 1;
  ram[27815]  = 1;
  ram[27816]  = 1;
  ram[27817]  = 1;
  ram[27818]  = 1;
  ram[27819]  = 1;
  ram[27820]  = 1;
  ram[27821]  = 1;
  ram[27822]  = 1;
  ram[27823]  = 1;
  ram[27824]  = 1;
  ram[27825]  = 1;
  ram[27826]  = 1;
  ram[27827]  = 1;
  ram[27828]  = 1;
  ram[27829]  = 1;
  ram[27830]  = 1;
  ram[27831]  = 1;
  ram[27832]  = 1;
  ram[27833]  = 1;
  ram[27834]  = 1;
  ram[27835]  = 1;
  ram[27836]  = 1;
  ram[27837]  = 1;
  ram[27838]  = 1;
  ram[27839]  = 1;
  ram[27840]  = 1;
  ram[27841]  = 1;
  ram[27842]  = 1;
  ram[27843]  = 1;
  ram[27844]  = 1;
  ram[27845]  = 1;
  ram[27846]  = 1;
  ram[27847]  = 1;
  ram[27848]  = 1;
  ram[27849]  = 1;
  ram[27850]  = 1;
  ram[27851]  = 1;
  ram[27852]  = 1;
  ram[27853]  = 1;
  ram[27854]  = 1;
  ram[27855]  = 1;
  ram[27856]  = 1;
  ram[27857]  = 1;
  ram[27858]  = 1;
  ram[27859]  = 1;
  ram[27860]  = 1;
  ram[27861]  = 1;
  ram[27862]  = 1;
  ram[27863]  = 1;
  ram[27864]  = 1;
  ram[27865]  = 1;
  ram[27866]  = 1;
  ram[27867]  = 1;
  ram[27868]  = 1;
  ram[27869]  = 1;
  ram[27870]  = 1;
  ram[27871]  = 1;
  ram[27872]  = 1;
  ram[27873]  = 1;
  ram[27874]  = 1;
  ram[27875]  = 1;
  ram[27876]  = 1;
  ram[27877]  = 1;
  ram[27878]  = 1;
  ram[27879]  = 1;
  ram[27880]  = 1;
  ram[27881]  = 1;
  ram[27882]  = 1;
  ram[27883]  = 1;
  ram[27884]  = 1;
  ram[27885]  = 1;
  ram[27886]  = 1;
  ram[27887]  = 1;
  ram[27888]  = 1;
  ram[27889]  = 1;
  ram[27890]  = 1;
  ram[27891]  = 1;
  ram[27892]  = 1;
  ram[27893]  = 1;
  ram[27894]  = 1;
  ram[27895]  = 1;
  ram[27896]  = 1;
  ram[27897]  = 1;
  ram[27898]  = 1;
  ram[27899]  = 1;
  ram[27900]  = 1;
  ram[27901]  = 1;
  ram[27902]  = 1;
  ram[27903]  = 1;
  ram[27904]  = 1;
  ram[27905]  = 1;
  ram[27906]  = 1;
  ram[27907]  = 1;
  ram[27908]  = 1;
  ram[27909]  = 1;
  ram[27910]  = 1;
  ram[27911]  = 1;
  ram[27912]  = 1;
  ram[27913]  = 1;
  ram[27914]  = 1;
  ram[27915]  = 1;
  ram[27916]  = 1;
  ram[27917]  = 1;
  ram[27918]  = 1;
  ram[27919]  = 1;
  ram[27920]  = 1;
  ram[27921]  = 1;
  ram[27922]  = 1;
  ram[27923]  = 1;
  ram[27924]  = 1;
  ram[27925]  = 1;
  ram[27926]  = 1;
  ram[27927]  = 1;
  ram[27928]  = 1;
  ram[27929]  = 1;
  ram[27930]  = 1;
  ram[27931]  = 1;
  ram[27932]  = 1;
  ram[27933]  = 1;
  ram[27934]  = 1;
  ram[27935]  = 1;
  ram[27936]  = 1;
  ram[27937]  = 1;
  ram[27938]  = 1;
  ram[27939]  = 1;
  ram[27940]  = 1;
  ram[27941]  = 1;
  ram[27942]  = 1;
  ram[27943]  = 1;
  ram[27944]  = 1;
  ram[27945]  = 1;
  ram[27946]  = 1;
  ram[27947]  = 1;
  ram[27948]  = 1;
  ram[27949]  = 1;
  ram[27950]  = 1;
  ram[27951]  = 1;
  ram[27952]  = 1;
  ram[27953]  = 1;
  ram[27954]  = 1;
  ram[27955]  = 1;
  ram[27956]  = 1;
  ram[27957]  = 1;
  ram[27958]  = 1;
  ram[27959]  = 1;
  ram[27960]  = 1;
  ram[27961]  = 1;
  ram[27962]  = 1;
  ram[27963]  = 1;
  ram[27964]  = 1;
  ram[27965]  = 1;
  ram[27966]  = 1;
  ram[27967]  = 1;
  ram[27968]  = 1;
  ram[27969]  = 1;
  ram[27970]  = 1;
  ram[27971]  = 1;
  ram[27972]  = 1;
  ram[27973]  = 1;
  ram[27974]  = 1;
  ram[27975]  = 1;
  ram[27976]  = 1;
  ram[27977]  = 1;
  ram[27978]  = 1;
  ram[27979]  = 1;
  ram[27980]  = 1;
  ram[27981]  = 1;
  ram[27982]  = 1;
  ram[27983]  = 1;
  ram[27984]  = 1;
  ram[27985]  = 1;
  ram[27986]  = 1;
  ram[27987]  = 1;
  ram[27988]  = 1;
  ram[27989]  = 1;
  ram[27990]  = 1;
  ram[27991]  = 1;
  ram[27992]  = 1;
  ram[27993]  = 1;
  ram[27994]  = 1;
  ram[27995]  = 1;
  ram[27996]  = 1;
  ram[27997]  = 1;
  ram[27998]  = 1;
  ram[27999]  = 1;
  ram[28000]  = 1;
  ram[28001]  = 1;
  ram[28002]  = 1;
  ram[28003]  = 1;
  ram[28004]  = 1;
  ram[28005]  = 1;
  ram[28006]  = 1;
  ram[28007]  = 1;
  ram[28008]  = 1;
  ram[28009]  = 1;
  ram[28010]  = 1;
  ram[28011]  = 1;
  ram[28012]  = 1;
  ram[28013]  = 1;
  ram[28014]  = 1;
  ram[28015]  = 1;
  ram[28016]  = 1;
  ram[28017]  = 1;
  ram[28018]  = 1;
  ram[28019]  = 1;
  ram[28020]  = 1;
  ram[28021]  = 1;
  ram[28022]  = 1;
  ram[28023]  = 1;
  ram[28024]  = 1;
  ram[28025]  = 1;
  ram[28026]  = 1;
  ram[28027]  = 1;
  ram[28028]  = 1;
  ram[28029]  = 1;
  ram[28030]  = 1;
  ram[28031]  = 1;
  ram[28032]  = 1;
  ram[28033]  = 1;
  ram[28034]  = 1;
  ram[28035]  = 1;
  ram[28036]  = 1;
  ram[28037]  = 1;
  ram[28038]  = 1;
  ram[28039]  = 1;
  ram[28040]  = 1;
  ram[28041]  = 1;
  ram[28042]  = 1;
  ram[28043]  = 1;
  ram[28044]  = 1;
  ram[28045]  = 1;
  ram[28046]  = 1;
  ram[28047]  = 1;
  ram[28048]  = 1;
  ram[28049]  = 1;
  ram[28050]  = 1;
  ram[28051]  = 1;
  ram[28052]  = 1;
  ram[28053]  = 1;
  ram[28054]  = 1;
  ram[28055]  = 1;
  ram[28056]  = 1;
  ram[28057]  = 1;
  ram[28058]  = 1;
  ram[28059]  = 1;
  ram[28060]  = 1;
  ram[28061]  = 1;
  ram[28062]  = 1;
  ram[28063]  = 1;
  ram[28064]  = 1;
  ram[28065]  = 1;
  ram[28066]  = 1;
  ram[28067]  = 1;
  ram[28068]  = 1;
  ram[28069]  = 1;
  ram[28070]  = 1;
  ram[28071]  = 1;
  ram[28072]  = 1;
  ram[28073]  = 1;
  ram[28074]  = 1;
  ram[28075]  = 1;
  ram[28076]  = 1;
  ram[28077]  = 1;
  ram[28078]  = 1;
  ram[28079]  = 1;
  ram[28080]  = 1;
  ram[28081]  = 1;
  ram[28082]  = 1;
  ram[28083]  = 1;
  ram[28084]  = 1;
  ram[28085]  = 1;
  ram[28086]  = 1;
  ram[28087]  = 1;
  ram[28088]  = 1;
  ram[28089]  = 1;
  ram[28090]  = 1;
  ram[28091]  = 1;
  ram[28092]  = 1;
  ram[28093]  = 1;
  ram[28094]  = 1;
  ram[28095]  = 1;
  ram[28096]  = 1;
  ram[28097]  = 1;
  ram[28098]  = 1;
  ram[28099]  = 1;
  ram[28100]  = 1;
  ram[28101]  = 1;
  ram[28102]  = 1;
  ram[28103]  = 1;
  ram[28104]  = 1;
  ram[28105]  = 1;
  ram[28106]  = 1;
  ram[28107]  = 1;
  ram[28108]  = 1;
  ram[28109]  = 1;
  ram[28110]  = 1;
  ram[28111]  = 1;
  ram[28112]  = 1;
  ram[28113]  = 1;
  ram[28114]  = 1;
  ram[28115]  = 1;
  ram[28116]  = 1;
  ram[28117]  = 1;
  ram[28118]  = 1;
  ram[28119]  = 1;
  ram[28120]  = 1;
  ram[28121]  = 1;
  ram[28122]  = 1;
  ram[28123]  = 1;
  ram[28124]  = 1;
  ram[28125]  = 1;
  ram[28126]  = 1;
  ram[28127]  = 1;
  ram[28128]  = 1;
  ram[28129]  = 1;
  ram[28130]  = 1;
  ram[28131]  = 1;
  ram[28132]  = 1;
  ram[28133]  = 1;
  ram[28134]  = 1;
  ram[28135]  = 1;
  ram[28136]  = 1;
  ram[28137]  = 1;
  ram[28138]  = 1;
  ram[28139]  = 1;
  ram[28140]  = 1;
  ram[28141]  = 1;
  ram[28142]  = 1;
  ram[28143]  = 1;
  ram[28144]  = 1;
  ram[28145]  = 1;
  ram[28146]  = 1;
  ram[28147]  = 1;
  ram[28148]  = 1;
  ram[28149]  = 1;
  ram[28150]  = 1;
  ram[28151]  = 1;
  ram[28152]  = 1;
  ram[28153]  = 1;
  ram[28154]  = 1;
  ram[28155]  = 1;
  ram[28156]  = 1;
  ram[28157]  = 1;
  ram[28158]  = 1;
  ram[28159]  = 1;
  ram[28160]  = 1;
  ram[28161]  = 1;
  ram[28162]  = 1;
  ram[28163]  = 1;
  ram[28164]  = 1;
  ram[28165]  = 1;
  ram[28166]  = 1;
  ram[28167]  = 1;
  ram[28168]  = 1;
  ram[28169]  = 1;
  ram[28170]  = 1;
  ram[28171]  = 1;
  ram[28172]  = 1;
  ram[28173]  = 1;
  ram[28174]  = 1;
  ram[28175]  = 1;
  ram[28176]  = 1;
  ram[28177]  = 1;
  ram[28178]  = 1;
  ram[28179]  = 1;
  ram[28180]  = 1;
  ram[28181]  = 1;
  ram[28182]  = 1;
  ram[28183]  = 1;
  ram[28184]  = 1;
  ram[28185]  = 1;
  ram[28186]  = 1;
  ram[28187]  = 1;
  ram[28188]  = 1;
  ram[28189]  = 1;
  ram[28190]  = 1;
  ram[28191]  = 1;
  ram[28192]  = 1;
  ram[28193]  = 1;
  ram[28194]  = 1;
  ram[28195]  = 1;
  ram[28196]  = 1;
  ram[28197]  = 1;
  ram[28198]  = 1;
  ram[28199]  = 1;
  ram[28200]  = 1;
  ram[28201]  = 1;
  ram[28202]  = 1;
  ram[28203]  = 1;
  ram[28204]  = 1;
  ram[28205]  = 1;
  ram[28206]  = 1;
  ram[28207]  = 1;
  ram[28208]  = 1;
  ram[28209]  = 1;
  ram[28210]  = 1;
  ram[28211]  = 1;
  ram[28212]  = 1;
  ram[28213]  = 1;
  ram[28214]  = 1;
  ram[28215]  = 1;
  ram[28216]  = 1;
  ram[28217]  = 1;
  ram[28218]  = 1;
  ram[28219]  = 1;
  ram[28220]  = 1;
  ram[28221]  = 1;
  ram[28222]  = 1;
  ram[28223]  = 1;
  ram[28224]  = 1;
  ram[28225]  = 1;
  ram[28226]  = 1;
  ram[28227]  = 1;
  ram[28228]  = 1;
  ram[28229]  = 1;
  ram[28230]  = 1;
  ram[28231]  = 1;
  ram[28232]  = 1;
  ram[28233]  = 1;
  ram[28234]  = 1;
  ram[28235]  = 1;
  ram[28236]  = 1;
  ram[28237]  = 1;
  ram[28238]  = 1;
  ram[28239]  = 1;
  ram[28240]  = 1;
  ram[28241]  = 1;
  ram[28242]  = 1;
  ram[28243]  = 1;
  ram[28244]  = 1;
  ram[28245]  = 1;
  ram[28246]  = 1;
  ram[28247]  = 1;
  ram[28248]  = 1;
  ram[28249]  = 1;
  ram[28250]  = 1;
  ram[28251]  = 1;
  ram[28252]  = 1;
  ram[28253]  = 1;
  ram[28254]  = 1;
  ram[28255]  = 1;
  ram[28256]  = 1;
  ram[28257]  = 1;
  ram[28258]  = 1;
  ram[28259]  = 1;
  ram[28260]  = 1;
  ram[28261]  = 1;
  ram[28262]  = 1;
  ram[28263]  = 1;
  ram[28264]  = 1;
  ram[28265]  = 1;
  ram[28266]  = 1;
  ram[28267]  = 1;
  ram[28268]  = 1;
  ram[28269]  = 1;
  ram[28270]  = 1;
  ram[28271]  = 1;
  ram[28272]  = 1;
  ram[28273]  = 1;
  ram[28274]  = 1;
  ram[28275]  = 1;
  ram[28276]  = 1;
  ram[28277]  = 1;
  ram[28278]  = 1;
  ram[28279]  = 1;
  ram[28280]  = 1;
  ram[28281]  = 1;
  ram[28282]  = 1;
  ram[28283]  = 1;
  ram[28284]  = 1;
  ram[28285]  = 1;
  ram[28286]  = 1;
  ram[28287]  = 1;
  ram[28288]  = 1;
  ram[28289]  = 1;
  ram[28290]  = 1;
  ram[28291]  = 1;
  ram[28292]  = 1;
  ram[28293]  = 1;
  ram[28294]  = 1;
  ram[28295]  = 1;
  ram[28296]  = 1;
  ram[28297]  = 1;
  ram[28298]  = 1;
  ram[28299]  = 1;
  ram[28300]  = 1;
  ram[28301]  = 1;
  ram[28302]  = 1;
  ram[28303]  = 1;
  ram[28304]  = 1;
  ram[28305]  = 1;
  ram[28306]  = 1;
  ram[28307]  = 1;
  ram[28308]  = 1;
  ram[28309]  = 1;
  ram[28310]  = 1;
  ram[28311]  = 1;
  ram[28312]  = 1;
  ram[28313]  = 1;
  ram[28314]  = 1;
  ram[28315]  = 1;
  ram[28316]  = 1;
  ram[28317]  = 1;
  ram[28318]  = 1;
  ram[28319]  = 1;
  ram[28320]  = 1;
  ram[28321]  = 1;
  ram[28322]  = 1;
  ram[28323]  = 1;
  ram[28324]  = 1;
  ram[28325]  = 1;
  ram[28326]  = 1;
  ram[28327]  = 1;
  ram[28328]  = 1;
  ram[28329]  = 1;
  ram[28330]  = 1;
  ram[28331]  = 1;
  ram[28332]  = 1;
  ram[28333]  = 1;
  ram[28334]  = 1;
  ram[28335]  = 1;
  ram[28336]  = 1;
  ram[28337]  = 1;
  ram[28338]  = 1;
  ram[28339]  = 1;
  ram[28340]  = 1;
  ram[28341]  = 1;
  ram[28342]  = 1;
  ram[28343]  = 1;
  ram[28344]  = 1;
  ram[28345]  = 1;
  ram[28346]  = 1;
  ram[28347]  = 1;
  ram[28348]  = 1;
  ram[28349]  = 1;
  ram[28350]  = 1;
  ram[28351]  = 1;
  ram[28352]  = 1;
  ram[28353]  = 1;
  ram[28354]  = 1;
  ram[28355]  = 1;
  ram[28356]  = 1;
  ram[28357]  = 1;
  ram[28358]  = 1;
  ram[28359]  = 1;
  ram[28360]  = 1;
  ram[28361]  = 1;
  ram[28362]  = 1;
  ram[28363]  = 1;
  ram[28364]  = 1;
  ram[28365]  = 1;
  ram[28366]  = 1;
  ram[28367]  = 1;
  ram[28368]  = 1;
  ram[28369]  = 1;
  ram[28370]  = 1;
  ram[28371]  = 1;
  ram[28372]  = 1;
  ram[28373]  = 1;
  ram[28374]  = 1;
  ram[28375]  = 1;
  ram[28376]  = 1;
  ram[28377]  = 1;
  ram[28378]  = 1;
  ram[28379]  = 1;
  ram[28380]  = 1;
  ram[28381]  = 1;
  ram[28382]  = 1;
  ram[28383]  = 1;
  ram[28384]  = 1;
  ram[28385]  = 1;
  ram[28386]  = 1;
  ram[28387]  = 1;
  ram[28388]  = 1;
  ram[28389]  = 1;
  ram[28390]  = 1;
  ram[28391]  = 1;
  ram[28392]  = 1;
  ram[28393]  = 1;
  ram[28394]  = 1;
  ram[28395]  = 1;
  ram[28396]  = 1;
  ram[28397]  = 1;
  ram[28398]  = 1;
  ram[28399]  = 1;
  ram[28400]  = 1;
  ram[28401]  = 1;
  ram[28402]  = 1;
  ram[28403]  = 1;
  ram[28404]  = 1;
  ram[28405]  = 1;
  ram[28406]  = 1;
  ram[28407]  = 1;
  ram[28408]  = 1;
  ram[28409]  = 1;
  ram[28410]  = 1;
  ram[28411]  = 1;
  ram[28412]  = 1;
  ram[28413]  = 1;
  ram[28414]  = 1;
  ram[28415]  = 1;
  ram[28416]  = 1;
  ram[28417]  = 1;
  ram[28418]  = 1;
  ram[28419]  = 1;
  ram[28420]  = 1;
  ram[28421]  = 1;
  ram[28422]  = 1;
  ram[28423]  = 1;
  ram[28424]  = 1;
  ram[28425]  = 1;
  ram[28426]  = 1;
  ram[28427]  = 1;
  ram[28428]  = 1;
  ram[28429]  = 1;
  ram[28430]  = 1;
  ram[28431]  = 1;
  ram[28432]  = 1;
  ram[28433]  = 1;
  ram[28434]  = 1;
  ram[28435]  = 1;
  ram[28436]  = 1;
  ram[28437]  = 1;
  ram[28438]  = 1;
  ram[28439]  = 1;
  ram[28440]  = 1;
  ram[28441]  = 1;
  ram[28442]  = 1;
  ram[28443]  = 1;
  ram[28444]  = 1;
  ram[28445]  = 1;
  ram[28446]  = 1;
  ram[28447]  = 1;
  ram[28448]  = 1;
  ram[28449]  = 1;
  ram[28450]  = 1;
  ram[28451]  = 1;
  ram[28452]  = 1;
  ram[28453]  = 1;
  ram[28454]  = 1;
  ram[28455]  = 1;
  ram[28456]  = 1;
  ram[28457]  = 1;
  ram[28458]  = 1;
  ram[28459]  = 1;
  ram[28460]  = 1;
  ram[28461]  = 1;
  ram[28462]  = 1;
  ram[28463]  = 1;
  ram[28464]  = 1;
  ram[28465]  = 1;
  ram[28466]  = 1;
  ram[28467]  = 1;
  ram[28468]  = 1;
  ram[28469]  = 1;
  ram[28470]  = 1;
  ram[28471]  = 1;
  ram[28472]  = 1;
  ram[28473]  = 1;
  ram[28474]  = 1;
  ram[28475]  = 1;
  ram[28476]  = 1;
  ram[28477]  = 1;
  ram[28478]  = 1;
  ram[28479]  = 1;
  ram[28480]  = 1;
  ram[28481]  = 1;
  ram[28482]  = 1;
  ram[28483]  = 1;
  ram[28484]  = 1;
  ram[28485]  = 1;
  ram[28486]  = 1;
  ram[28487]  = 1;
  ram[28488]  = 1;
  ram[28489]  = 1;
  ram[28490]  = 1;
  ram[28491]  = 1;
  ram[28492]  = 1;
  ram[28493]  = 1;
  ram[28494]  = 1;
  ram[28495]  = 1;
  ram[28496]  = 1;
  ram[28497]  = 1;
  ram[28498]  = 1;
  ram[28499]  = 1;
  ram[28500]  = 1;
  ram[28501]  = 1;
  ram[28502]  = 1;
  ram[28503]  = 1;
  ram[28504]  = 1;
  ram[28505]  = 1;
  ram[28506]  = 1;
  ram[28507]  = 1;
  ram[28508]  = 1;
  ram[28509]  = 1;
  ram[28510]  = 1;
  ram[28511]  = 1;
  ram[28512]  = 1;
  ram[28513]  = 1;
  ram[28514]  = 1;
  ram[28515]  = 1;
  ram[28516]  = 1;
  ram[28517]  = 1;
  ram[28518]  = 1;
  ram[28519]  = 1;
  ram[28520]  = 1;
  ram[28521]  = 1;
  ram[28522]  = 1;
  ram[28523]  = 1;
  ram[28524]  = 1;
  ram[28525]  = 1;
  ram[28526]  = 1;
  ram[28527]  = 1;
  ram[28528]  = 1;
  ram[28529]  = 1;
  ram[28530]  = 1;
  ram[28531]  = 1;
  ram[28532]  = 1;
  ram[28533]  = 1;
  ram[28534]  = 1;
  ram[28535]  = 1;
  ram[28536]  = 1;
  ram[28537]  = 1;
  ram[28538]  = 1;
  ram[28539]  = 1;
  ram[28540]  = 1;
  ram[28541]  = 1;
  ram[28542]  = 1;
  ram[28543]  = 1;
  ram[28544]  = 1;
  ram[28545]  = 1;
  ram[28546]  = 1;
  ram[28547]  = 1;
  ram[28548]  = 1;
  ram[28549]  = 1;
  ram[28550]  = 1;
  ram[28551]  = 1;
  ram[28552]  = 1;
  ram[28553]  = 1;
  ram[28554]  = 1;
  ram[28555]  = 1;
  ram[28556]  = 1;
  ram[28557]  = 1;
  ram[28558]  = 1;
  ram[28559]  = 1;
  ram[28560]  = 1;
  ram[28561]  = 1;
  ram[28562]  = 1;
  ram[28563]  = 1;
  ram[28564]  = 1;
  ram[28565]  = 1;
  ram[28566]  = 1;
  ram[28567]  = 1;
  ram[28568]  = 1;
  ram[28569]  = 1;
  ram[28570]  = 1;
  ram[28571]  = 1;
  ram[28572]  = 1;
  ram[28573]  = 1;
  ram[28574]  = 1;
  ram[28575]  = 1;
  ram[28576]  = 1;
  ram[28577]  = 1;
  ram[28578]  = 1;
  ram[28579]  = 1;
  ram[28580]  = 1;
  ram[28581]  = 1;
  ram[28582]  = 1;
  ram[28583]  = 1;
  ram[28584]  = 1;
  ram[28585]  = 1;
  ram[28586]  = 1;
  ram[28587]  = 1;
  ram[28588]  = 1;
  ram[28589]  = 1;
  ram[28590]  = 1;
  ram[28591]  = 1;
  ram[28592]  = 1;
  ram[28593]  = 1;
  ram[28594]  = 1;
  ram[28595]  = 1;
  ram[28596]  = 1;
  ram[28597]  = 1;
  ram[28598]  = 1;
  ram[28599]  = 1;
  ram[28600]  = 1;
  ram[28601]  = 1;
  ram[28602]  = 1;
  ram[28603]  = 1;
  ram[28604]  = 1;
  ram[28605]  = 1;
  ram[28606]  = 1;
  ram[28607]  = 1;
  ram[28608]  = 1;
  ram[28609]  = 1;
  ram[28610]  = 1;
  ram[28611]  = 1;
  ram[28612]  = 1;
  ram[28613]  = 1;
  ram[28614]  = 1;
  ram[28615]  = 1;
  ram[28616]  = 1;
  ram[28617]  = 1;
  ram[28618]  = 1;
  ram[28619]  = 1;
  ram[28620]  = 1;
  ram[28621]  = 1;
  ram[28622]  = 1;
  ram[28623]  = 1;
  ram[28624]  = 1;
  ram[28625]  = 1;
  ram[28626]  = 1;
  ram[28627]  = 1;
  ram[28628]  = 1;
  ram[28629]  = 1;
  ram[28630]  = 1;
  ram[28631]  = 1;
  ram[28632]  = 1;
  ram[28633]  = 1;
  ram[28634]  = 1;
  ram[28635]  = 1;
  ram[28636]  = 1;
  ram[28637]  = 1;
  ram[28638]  = 1;
  ram[28639]  = 1;
  ram[28640]  = 1;
  ram[28641]  = 1;
  ram[28642]  = 1;
  ram[28643]  = 1;
  ram[28644]  = 1;
  ram[28645]  = 1;
  ram[28646]  = 1;
  ram[28647]  = 1;
  ram[28648]  = 1;
  ram[28649]  = 1;
  ram[28650]  = 1;
  ram[28651]  = 1;
  ram[28652]  = 1;
  ram[28653]  = 1;
  ram[28654]  = 1;
  ram[28655]  = 1;
  ram[28656]  = 1;
  ram[28657]  = 1;
  ram[28658]  = 1;
  ram[28659]  = 1;
  ram[28660]  = 1;
  ram[28661]  = 1;
  ram[28662]  = 1;
  ram[28663]  = 1;
  ram[28664]  = 1;
  ram[28665]  = 1;
  ram[28666]  = 1;
  ram[28667]  = 1;
  ram[28668]  = 1;
  ram[28669]  = 1;
  ram[28670]  = 1;
  ram[28671]  = 1;
  ram[28672]  = 1;
  ram[28673]  = 1;
  ram[28674]  = 1;
  ram[28675]  = 1;
  ram[28676]  = 1;
  ram[28677]  = 1;
  ram[28678]  = 1;
  ram[28679]  = 1;
  ram[28680]  = 1;
  ram[28681]  = 1;
  ram[28682]  = 1;
  ram[28683]  = 1;
  ram[28684]  = 1;
  ram[28685]  = 1;
  ram[28686]  = 1;
  ram[28687]  = 1;
  ram[28688]  = 1;
  ram[28689]  = 1;
  ram[28690]  = 1;
  ram[28691]  = 1;
  ram[28692]  = 1;
  ram[28693]  = 1;
  ram[28694]  = 1;
  ram[28695]  = 1;
  ram[28696]  = 1;
  ram[28697]  = 1;
  ram[28698]  = 1;
  ram[28699]  = 1;
  ram[28700]  = 1;
  ram[28701]  = 1;
  ram[28702]  = 1;
  ram[28703]  = 1;
  ram[28704]  = 1;
  ram[28705]  = 1;
  ram[28706]  = 1;
  ram[28707]  = 1;
  ram[28708]  = 1;
  ram[28709]  = 1;
  ram[28710]  = 1;
  ram[28711]  = 1;
  ram[28712]  = 1;
  ram[28713]  = 1;
  ram[28714]  = 1;
  ram[28715]  = 1;
  ram[28716]  = 1;
  ram[28717]  = 1;
  ram[28718]  = 1;
  ram[28719]  = 1;
  ram[28720]  = 1;
  ram[28721]  = 1;
  ram[28722]  = 1;
  ram[28723]  = 1;
  ram[28724]  = 1;
  ram[28725]  = 1;
  ram[28726]  = 1;
  ram[28727]  = 1;
  ram[28728]  = 1;
  ram[28729]  = 1;
  ram[28730]  = 1;
  ram[28731]  = 1;
  ram[28732]  = 1;
  ram[28733]  = 1;
  ram[28734]  = 1;
  ram[28735]  = 1;
  ram[28736]  = 1;
  ram[28737]  = 1;
  ram[28738]  = 1;
  ram[28739]  = 1;
  ram[28740]  = 1;
  ram[28741]  = 1;
  ram[28742]  = 1;
  ram[28743]  = 1;
  ram[28744]  = 1;
  ram[28745]  = 1;
  ram[28746]  = 1;
  ram[28747]  = 1;
  ram[28748]  = 1;
  ram[28749]  = 1;
  ram[28750]  = 1;
  ram[28751]  = 1;
  ram[28752]  = 1;
  ram[28753]  = 1;
  ram[28754]  = 1;
  ram[28755]  = 1;
  ram[28756]  = 1;
  ram[28757]  = 1;
  ram[28758]  = 1;
  ram[28759]  = 1;
  ram[28760]  = 1;
  ram[28761]  = 1;
  ram[28762]  = 1;
  ram[28763]  = 1;
  ram[28764]  = 1;
  ram[28765]  = 1;
  ram[28766]  = 1;
  ram[28767]  = 1;
  ram[28768]  = 1;
  ram[28769]  = 1;
  ram[28770]  = 1;
  ram[28771]  = 1;
  ram[28772]  = 1;
  ram[28773]  = 1;
  ram[28774]  = 1;
  ram[28775]  = 1;
  ram[28776]  = 1;
  ram[28777]  = 1;
  ram[28778]  = 1;
  ram[28779]  = 1;
  ram[28780]  = 1;
  ram[28781]  = 1;
  ram[28782]  = 1;
  ram[28783]  = 1;
  ram[28784]  = 1;
  ram[28785]  = 1;
  ram[28786]  = 1;
  ram[28787]  = 1;
  ram[28788]  = 1;
  ram[28789]  = 1;
  ram[28790]  = 1;
  ram[28791]  = 1;
  ram[28792]  = 1;
  ram[28793]  = 1;
  ram[28794]  = 1;
  ram[28795]  = 1;
  ram[28796]  = 1;
  ram[28797]  = 1;
  ram[28798]  = 1;
  ram[28799]  = 1;
  ram[28800]  = 1;
  ram[28801]  = 1;
  ram[28802]  = 1;
  ram[28803]  = 1;
  ram[28804]  = 1;
  ram[28805]  = 1;
  ram[28806]  = 1;
  ram[28807]  = 1;
  ram[28808]  = 1;
  ram[28809]  = 1;
  ram[28810]  = 1;
  ram[28811]  = 1;
  ram[28812]  = 1;
  ram[28813]  = 1;
  ram[28814]  = 1;
  ram[28815]  = 1;
  ram[28816]  = 1;
  ram[28817]  = 1;
  ram[28818]  = 1;
  ram[28819]  = 1;
  ram[28820]  = 1;
  ram[28821]  = 1;
  ram[28822]  = 1;
  ram[28823]  = 1;
  ram[28824]  = 1;
  ram[28825]  = 1;
  ram[28826]  = 1;
  ram[28827]  = 1;
  ram[28828]  = 1;
  ram[28829]  = 1;
  ram[28830]  = 1;
  ram[28831]  = 1;
  ram[28832]  = 1;
  ram[28833]  = 1;
  ram[28834]  = 1;
  ram[28835]  = 1;
  ram[28836]  = 1;
  ram[28837]  = 1;
  ram[28838]  = 1;
  ram[28839]  = 1;
  ram[28840]  = 1;
  ram[28841]  = 1;
  ram[28842]  = 1;
  ram[28843]  = 1;
  ram[28844]  = 1;
  ram[28845]  = 1;
  ram[28846]  = 1;
  ram[28847]  = 1;
  ram[28848]  = 1;
  ram[28849]  = 1;
  ram[28850]  = 1;
  ram[28851]  = 1;
  ram[28852]  = 1;
  ram[28853]  = 1;
  ram[28854]  = 1;
  ram[28855]  = 1;
  ram[28856]  = 1;
  ram[28857]  = 1;
  ram[28858]  = 1;
  ram[28859]  = 1;
  ram[28860]  = 1;
  ram[28861]  = 1;
  ram[28862]  = 1;
  ram[28863]  = 1;
  ram[28864]  = 1;
  ram[28865]  = 1;
  ram[28866]  = 1;
  ram[28867]  = 1;
  ram[28868]  = 1;
  ram[28869]  = 1;
  ram[28870]  = 1;
  ram[28871]  = 1;
  ram[28872]  = 1;
  ram[28873]  = 1;
  ram[28874]  = 1;
  ram[28875]  = 1;
  ram[28876]  = 1;
  ram[28877]  = 1;
  ram[28878]  = 1;
  ram[28879]  = 1;
  ram[28880]  = 1;
  ram[28881]  = 1;
  ram[28882]  = 1;
  ram[28883]  = 1;
  ram[28884]  = 1;
  ram[28885]  = 1;
  ram[28886]  = 1;
  ram[28887]  = 1;
  ram[28888]  = 1;
  ram[28889]  = 1;
  ram[28890]  = 1;
  ram[28891]  = 1;
  ram[28892]  = 1;
  ram[28893]  = 1;
  ram[28894]  = 1;
  ram[28895]  = 1;
  ram[28896]  = 1;
  ram[28897]  = 1;
  ram[28898]  = 1;
  ram[28899]  = 1;
  ram[28900]  = 1;
  ram[28901]  = 1;
  ram[28902]  = 1;
  ram[28903]  = 1;
  ram[28904]  = 1;
  ram[28905]  = 1;
  ram[28906]  = 1;
  ram[28907]  = 1;
  ram[28908]  = 1;
  ram[28909]  = 1;
  ram[28910]  = 1;
  ram[28911]  = 1;
  ram[28912]  = 1;
  ram[28913]  = 1;
  ram[28914]  = 1;
  ram[28915]  = 1;
  ram[28916]  = 1;
  ram[28917]  = 1;
  ram[28918]  = 1;
  ram[28919]  = 1;
  ram[28920]  = 1;
  ram[28921]  = 1;
  ram[28922]  = 1;
  ram[28923]  = 1;
  ram[28924]  = 1;
  ram[28925]  = 1;
  ram[28926]  = 1;
  ram[28927]  = 1;
  ram[28928]  = 1;
  ram[28929]  = 1;
  ram[28930]  = 1;
  ram[28931]  = 1;
  ram[28932]  = 1;
  ram[28933]  = 1;
  ram[28934]  = 1;
  ram[28935]  = 1;
  ram[28936]  = 1;
  ram[28937]  = 1;
  ram[28938]  = 1;
  ram[28939]  = 1;
  ram[28940]  = 1;
  ram[28941]  = 1;
  ram[28942]  = 1;
  ram[28943]  = 1;
  ram[28944]  = 1;
  ram[28945]  = 1;
  ram[28946]  = 1;
  ram[28947]  = 1;
  ram[28948]  = 1;
  ram[28949]  = 1;
  ram[28950]  = 1;
  ram[28951]  = 1;
  ram[28952]  = 1;
  ram[28953]  = 1;
  ram[28954]  = 1;
  ram[28955]  = 1;
  ram[28956]  = 1;
  ram[28957]  = 1;
  ram[28958]  = 1;
  ram[28959]  = 1;
  ram[28960]  = 1;
  ram[28961]  = 1;
  ram[28962]  = 1;
  ram[28963]  = 1;
  ram[28964]  = 1;
  ram[28965]  = 1;
  ram[28966]  = 1;
  ram[28967]  = 1;
  ram[28968]  = 1;
  ram[28969]  = 1;
  ram[28970]  = 1;
  ram[28971]  = 1;
  ram[28972]  = 1;
  ram[28973]  = 1;
  ram[28974]  = 1;
  ram[28975]  = 1;
  ram[28976]  = 1;
  ram[28977]  = 1;
  ram[28978]  = 1;
  ram[28979]  = 1;
  ram[28980]  = 1;
  ram[28981]  = 1;
  ram[28982]  = 1;
  ram[28983]  = 1;
  ram[28984]  = 1;
  ram[28985]  = 1;
  ram[28986]  = 1;
  ram[28987]  = 1;
  ram[28988]  = 1;
  ram[28989]  = 1;
  ram[28990]  = 1;
  ram[28991]  = 1;
  ram[28992]  = 1;
  ram[28993]  = 1;
  ram[28994]  = 1;
  ram[28995]  = 1;
  ram[28996]  = 1;
  ram[28997]  = 1;
  ram[28998]  = 1;
  ram[28999]  = 1;
  ram[29000]  = 1;
  ram[29001]  = 1;
  ram[29002]  = 1;
  ram[29003]  = 1;
  ram[29004]  = 1;
  ram[29005]  = 1;
  ram[29006]  = 1;
  ram[29007]  = 1;
  ram[29008]  = 1;
  ram[29009]  = 1;
  ram[29010]  = 1;
  ram[29011]  = 1;
  ram[29012]  = 1;
  ram[29013]  = 1;
  ram[29014]  = 1;
  ram[29015]  = 1;
  ram[29016]  = 1;
  ram[29017]  = 1;
  ram[29018]  = 1;
  ram[29019]  = 1;
  ram[29020]  = 1;
  ram[29021]  = 1;
  ram[29022]  = 1;
  ram[29023]  = 1;
  ram[29024]  = 1;
  ram[29025]  = 1;
  ram[29026]  = 1;
  ram[29027]  = 1;
  ram[29028]  = 1;
  ram[29029]  = 1;
  ram[29030]  = 1;
  ram[29031]  = 1;
  ram[29032]  = 1;
  ram[29033]  = 1;
  ram[29034]  = 1;
  ram[29035]  = 1;
  ram[29036]  = 1;
  ram[29037]  = 1;
  ram[29038]  = 1;
  ram[29039]  = 1;
  ram[29040]  = 1;
  ram[29041]  = 1;
  ram[29042]  = 1;
  ram[29043]  = 1;
  ram[29044]  = 1;
  ram[29045]  = 1;
  ram[29046]  = 1;
  ram[29047]  = 1;
  ram[29048]  = 1;
  ram[29049]  = 1;
  ram[29050]  = 1;
  ram[29051]  = 1;
  ram[29052]  = 1;
  ram[29053]  = 1;
  ram[29054]  = 1;
  ram[29055]  = 1;
  ram[29056]  = 1;
  ram[29057]  = 1;
  ram[29058]  = 1;
  ram[29059]  = 1;
  ram[29060]  = 1;
  ram[29061]  = 1;
  ram[29062]  = 1;
  ram[29063]  = 1;
  ram[29064]  = 1;
  ram[29065]  = 1;
  ram[29066]  = 1;
  ram[29067]  = 1;
  ram[29068]  = 1;
  ram[29069]  = 1;
  ram[29070]  = 1;
  ram[29071]  = 1;
  ram[29072]  = 1;
  ram[29073]  = 1;
  ram[29074]  = 1;
  ram[29075]  = 1;
  ram[29076]  = 1;
  ram[29077]  = 1;
  ram[29078]  = 1;
  ram[29079]  = 1;
  ram[29080]  = 1;
  ram[29081]  = 1;
  ram[29082]  = 1;
  ram[29083]  = 1;
  ram[29084]  = 1;
  ram[29085]  = 1;
  ram[29086]  = 1;
  ram[29087]  = 1;
  ram[29088]  = 1;
  ram[29089]  = 1;
  ram[29090]  = 1;
  ram[29091]  = 1;
  ram[29092]  = 1;
  ram[29093]  = 1;
  ram[29094]  = 1;
  ram[29095]  = 1;
  ram[29096]  = 1;
  ram[29097]  = 1;
  ram[29098]  = 1;
  ram[29099]  = 1;
  ram[29100]  = 1;
  ram[29101]  = 1;
  ram[29102]  = 1;
  ram[29103]  = 1;
  ram[29104]  = 1;
  ram[29105]  = 1;
  ram[29106]  = 1;
  ram[29107]  = 1;
  ram[29108]  = 1;
  ram[29109]  = 1;
  ram[29110]  = 1;
  ram[29111]  = 1;
  ram[29112]  = 1;
  ram[29113]  = 1;
  ram[29114]  = 1;
  ram[29115]  = 1;
  ram[29116]  = 1;
  ram[29117]  = 1;
  ram[29118]  = 1;
  ram[29119]  = 1;
  ram[29120]  = 1;
  ram[29121]  = 1;
  ram[29122]  = 1;
  ram[29123]  = 1;
  ram[29124]  = 1;
  ram[29125]  = 1;
  ram[29126]  = 1;
  ram[29127]  = 1;
  ram[29128]  = 1;
  ram[29129]  = 1;
  ram[29130]  = 1;
  ram[29131]  = 1;
  ram[29132]  = 1;
  ram[29133]  = 1;
  ram[29134]  = 1;
  ram[29135]  = 1;
  ram[29136]  = 1;
  ram[29137]  = 1;
  ram[29138]  = 1;
  ram[29139]  = 1;
  ram[29140]  = 1;
  ram[29141]  = 1;
  ram[29142]  = 1;
  ram[29143]  = 1;
  ram[29144]  = 1;
  ram[29145]  = 1;
  ram[29146]  = 1;
  ram[29147]  = 1;
  ram[29148]  = 1;
  ram[29149]  = 1;
  ram[29150]  = 1;
  ram[29151]  = 1;
  ram[29152]  = 1;
  ram[29153]  = 1;
  ram[29154]  = 1;
  ram[29155]  = 1;
  ram[29156]  = 1;
  ram[29157]  = 1;
  ram[29158]  = 1;
  ram[29159]  = 1;
  ram[29160]  = 1;
  ram[29161]  = 1;
  ram[29162]  = 1;
  ram[29163]  = 1;
  ram[29164]  = 1;
  ram[29165]  = 1;
  ram[29166]  = 1;
  ram[29167]  = 1;
  ram[29168]  = 1;
  ram[29169]  = 1;
  ram[29170]  = 1;
  ram[29171]  = 1;
  ram[29172]  = 1;
  ram[29173]  = 1;
  ram[29174]  = 1;
  ram[29175]  = 1;
  ram[29176]  = 1;
  ram[29177]  = 1;
  ram[29178]  = 1;
  ram[29179]  = 1;
  ram[29180]  = 1;
  ram[29181]  = 1;
  ram[29182]  = 1;
  ram[29183]  = 1;
  ram[29184]  = 1;
  ram[29185]  = 1;
  ram[29186]  = 1;
  ram[29187]  = 1;
  ram[29188]  = 1;
  ram[29189]  = 1;
  ram[29190]  = 1;
  ram[29191]  = 1;
  ram[29192]  = 1;
  ram[29193]  = 1;
  ram[29194]  = 1;
  ram[29195]  = 1;
  ram[29196]  = 1;
  ram[29197]  = 1;
  ram[29198]  = 1;
  ram[29199]  = 1;
  ram[29200]  = 1;
  ram[29201]  = 1;
  ram[29202]  = 1;
  ram[29203]  = 1;
  ram[29204]  = 1;
  ram[29205]  = 1;
  ram[29206]  = 1;
  ram[29207]  = 1;
  ram[29208]  = 1;
  ram[29209]  = 1;
  ram[29210]  = 1;
  ram[29211]  = 1;
  ram[29212]  = 1;
  ram[29213]  = 1;
  ram[29214]  = 1;
  ram[29215]  = 1;
  ram[29216]  = 1;
  ram[29217]  = 1;
  ram[29218]  = 1;
  ram[29219]  = 1;
  ram[29220]  = 1;
  ram[29221]  = 1;
  ram[29222]  = 1;
  ram[29223]  = 1;
  ram[29224]  = 1;
  ram[29225]  = 1;
  ram[29226]  = 1;
  ram[29227]  = 1;
  ram[29228]  = 1;
  ram[29229]  = 1;
  ram[29230]  = 1;
  ram[29231]  = 1;
  ram[29232]  = 1;
  ram[29233]  = 1;
  ram[29234]  = 1;
  ram[29235]  = 1;
  ram[29236]  = 1;
  ram[29237]  = 1;
  ram[29238]  = 1;
  ram[29239]  = 1;
  ram[29240]  = 1;
  ram[29241]  = 1;
  ram[29242]  = 1;
  ram[29243]  = 1;
  ram[29244]  = 1;
  ram[29245]  = 1;
  ram[29246]  = 1;
  ram[29247]  = 1;
  ram[29248]  = 1;
  ram[29249]  = 1;
  ram[29250]  = 1;
  ram[29251]  = 1;
  ram[29252]  = 1;
  ram[29253]  = 1;
  ram[29254]  = 1;
  ram[29255]  = 1;
  ram[29256]  = 1;
  ram[29257]  = 1;
  ram[29258]  = 1;
  ram[29259]  = 1;
  ram[29260]  = 1;
  ram[29261]  = 1;
  ram[29262]  = 1;
  ram[29263]  = 1;
  ram[29264]  = 1;
  ram[29265]  = 1;
  ram[29266]  = 1;
  ram[29267]  = 1;
  ram[29268]  = 1;
  ram[29269]  = 1;
  ram[29270]  = 1;
  ram[29271]  = 1;
  ram[29272]  = 1;
  ram[29273]  = 1;
  ram[29274]  = 1;
  ram[29275]  = 1;
  ram[29276]  = 1;
  ram[29277]  = 1;
  ram[29278]  = 1;
  ram[29279]  = 1;
  ram[29280]  = 1;
  ram[29281]  = 1;
  ram[29282]  = 1;
  ram[29283]  = 1;
  ram[29284]  = 1;
  ram[29285]  = 1;
  ram[29286]  = 1;
  ram[29287]  = 1;
  ram[29288]  = 1;
  ram[29289]  = 1;
  ram[29290]  = 1;
  ram[29291]  = 1;
  ram[29292]  = 1;
  ram[29293]  = 1;
  ram[29294]  = 1;
  ram[29295]  = 1;
  ram[29296]  = 1;
  ram[29297]  = 1;
  ram[29298]  = 1;
  ram[29299]  = 1;
  ram[29300]  = 1;
  ram[29301]  = 1;
  ram[29302]  = 1;
  ram[29303]  = 1;
  ram[29304]  = 1;
  ram[29305]  = 1;
  ram[29306]  = 1;
  ram[29307]  = 1;
  ram[29308]  = 1;
  ram[29309]  = 1;
  ram[29310]  = 1;
  ram[29311]  = 1;
  ram[29312]  = 1;
  ram[29313]  = 1;
  ram[29314]  = 1;
  ram[29315]  = 1;
  ram[29316]  = 1;
  ram[29317]  = 1;
  ram[29318]  = 1;
  ram[29319]  = 1;
  ram[29320]  = 1;
  ram[29321]  = 1;
  ram[29322]  = 1;
  ram[29323]  = 1;
  ram[29324]  = 1;
  ram[29325]  = 1;
  ram[29326]  = 1;
  ram[29327]  = 1;
  ram[29328]  = 1;
  ram[29329]  = 1;
  ram[29330]  = 1;
  ram[29331]  = 1;
  ram[29332]  = 1;
  ram[29333]  = 1;
  ram[29334]  = 1;
  ram[29335]  = 1;
  ram[29336]  = 1;
  ram[29337]  = 1;
  ram[29338]  = 1;
  ram[29339]  = 1;
  ram[29340]  = 1;
  ram[29341]  = 1;
  ram[29342]  = 1;
  ram[29343]  = 1;
  ram[29344]  = 1;
  ram[29345]  = 1;
  ram[29346]  = 1;
  ram[29347]  = 1;
  ram[29348]  = 1;
  ram[29349]  = 1;
  ram[29350]  = 1;
  ram[29351]  = 1;
  ram[29352]  = 1;
  ram[29353]  = 1;
  ram[29354]  = 1;
  ram[29355]  = 1;
  ram[29356]  = 1;
  ram[29357]  = 1;
  ram[29358]  = 1;
  ram[29359]  = 1;
  ram[29360]  = 1;
  ram[29361]  = 1;
  ram[29362]  = 1;
  ram[29363]  = 1;
  ram[29364]  = 1;
  ram[29365]  = 1;
  ram[29366]  = 1;
  ram[29367]  = 1;
  ram[29368]  = 1;
  ram[29369]  = 1;
  ram[29370]  = 1;
  ram[29371]  = 1;
  ram[29372]  = 1;
  ram[29373]  = 1;
  ram[29374]  = 1;
  ram[29375]  = 1;
  ram[29376]  = 1;
  ram[29377]  = 1;
  ram[29378]  = 1;
  ram[29379]  = 1;
  ram[29380]  = 1;
  ram[29381]  = 1;
  ram[29382]  = 1;
  ram[29383]  = 1;
  ram[29384]  = 1;
  ram[29385]  = 1;
  ram[29386]  = 1;
  ram[29387]  = 1;
  ram[29388]  = 1;
  ram[29389]  = 1;
  ram[29390]  = 1;
  ram[29391]  = 1;
  ram[29392]  = 1;
  ram[29393]  = 1;
  ram[29394]  = 1;
  ram[29395]  = 1;
  ram[29396]  = 1;
  ram[29397]  = 1;
  ram[29398]  = 1;
  ram[29399]  = 1;
  ram[29400]  = 1;
  ram[29401]  = 1;
  ram[29402]  = 1;
  ram[29403]  = 1;
  ram[29404]  = 1;
  ram[29405]  = 1;
  ram[29406]  = 1;
  ram[29407]  = 1;
  ram[29408]  = 1;
  ram[29409]  = 1;
  ram[29410]  = 1;
  ram[29411]  = 1;
  ram[29412]  = 1;
  ram[29413]  = 1;
  ram[29414]  = 1;
  ram[29415]  = 1;
  ram[29416]  = 1;
  ram[29417]  = 1;
  ram[29418]  = 1;
  ram[29419]  = 1;
  ram[29420]  = 1;
  ram[29421]  = 1;
  ram[29422]  = 1;
  ram[29423]  = 1;
  ram[29424]  = 1;
  ram[29425]  = 1;
  ram[29426]  = 1;
  ram[29427]  = 1;
  ram[29428]  = 1;
  ram[29429]  = 1;
  ram[29430]  = 1;
  ram[29431]  = 1;
  ram[29432]  = 1;
  ram[29433]  = 1;
  ram[29434]  = 1;
  ram[29435]  = 1;
  ram[29436]  = 1;
  ram[29437]  = 1;
  ram[29438]  = 1;
  ram[29439]  = 1;
  ram[29440]  = 1;
  ram[29441]  = 1;
  ram[29442]  = 1;
  ram[29443]  = 1;
  ram[29444]  = 1;
  ram[29445]  = 1;
  ram[29446]  = 1;
  ram[29447]  = 1;
  ram[29448]  = 1;
  ram[29449]  = 1;
  ram[29450]  = 1;
  ram[29451]  = 1;
  ram[29452]  = 1;
  ram[29453]  = 1;
  ram[29454]  = 1;
  ram[29455]  = 1;
  ram[29456]  = 1;
  ram[29457]  = 1;
  ram[29458]  = 1;
  ram[29459]  = 1;
  ram[29460]  = 1;
  ram[29461]  = 1;
  ram[29462]  = 1;
  ram[29463]  = 1;
  ram[29464]  = 1;
  ram[29465]  = 1;
  ram[29466]  = 1;
  ram[29467]  = 1;
  ram[29468]  = 1;
  ram[29469]  = 1;
  ram[29470]  = 1;
  ram[29471]  = 1;
  ram[29472]  = 1;
  ram[29473]  = 1;
  ram[29474]  = 1;
  ram[29475]  = 1;
  ram[29476]  = 1;
  ram[29477]  = 1;
  ram[29478]  = 1;
  ram[29479]  = 1;
  ram[29480]  = 1;
  ram[29481]  = 1;
  ram[29482]  = 1;
  ram[29483]  = 1;
  ram[29484]  = 1;
  ram[29485]  = 1;
  ram[29486]  = 1;
  ram[29487]  = 1;
  ram[29488]  = 1;
  ram[29489]  = 1;
  ram[29490]  = 1;
  ram[29491]  = 1;
  ram[29492]  = 1;
  ram[29493]  = 1;
  ram[29494]  = 1;
  ram[29495]  = 1;
  ram[29496]  = 1;
  ram[29497]  = 1;
  ram[29498]  = 1;
  ram[29499]  = 1;
  ram[29500]  = 1;
  ram[29501]  = 1;
  ram[29502]  = 1;
  ram[29503]  = 1;
  ram[29504]  = 1;
  ram[29505]  = 1;
  ram[29506]  = 1;
  ram[29507]  = 1;
  ram[29508]  = 1;
  ram[29509]  = 1;
  ram[29510]  = 1;
  ram[29511]  = 1;
  ram[29512]  = 1;
  ram[29513]  = 1;
  ram[29514]  = 1;
  ram[29515]  = 1;
  ram[29516]  = 1;
  ram[29517]  = 1;
  ram[29518]  = 1;
  ram[29519]  = 1;
  ram[29520]  = 1;
  ram[29521]  = 1;
  ram[29522]  = 1;
  ram[29523]  = 1;
  ram[29524]  = 1;
  ram[29525]  = 1;
  ram[29526]  = 1;
  ram[29527]  = 1;
  ram[29528]  = 1;
  ram[29529]  = 1;
  ram[29530]  = 1;
  ram[29531]  = 1;
  ram[29532]  = 1;
  ram[29533]  = 1;
  ram[29534]  = 1;
  ram[29535]  = 1;
  ram[29536]  = 1;
  ram[29537]  = 1;
  ram[29538]  = 1;
  ram[29539]  = 1;
  ram[29540]  = 1;
  ram[29541]  = 1;
  ram[29542]  = 1;
  ram[29543]  = 1;
  ram[29544]  = 1;
  ram[29545]  = 1;
  ram[29546]  = 1;
  ram[29547]  = 1;
  ram[29548]  = 1;
  ram[29549]  = 1;
  ram[29550]  = 1;
  ram[29551]  = 1;
  ram[29552]  = 1;
  ram[29553]  = 1;
  ram[29554]  = 1;
  ram[29555]  = 1;
  ram[29556]  = 1;
  ram[29557]  = 1;
  ram[29558]  = 1;
  ram[29559]  = 1;
  ram[29560]  = 1;
  ram[29561]  = 1;
  ram[29562]  = 1;
  ram[29563]  = 1;
  ram[29564]  = 1;
  ram[29565]  = 1;
  ram[29566]  = 1;
  ram[29567]  = 1;
  ram[29568]  = 1;
  ram[29569]  = 1;
  ram[29570]  = 1;
  ram[29571]  = 1;
  ram[29572]  = 1;
  ram[29573]  = 1;
  ram[29574]  = 1;
  ram[29575]  = 1;
  ram[29576]  = 1;
  ram[29577]  = 1;
  ram[29578]  = 1;
  ram[29579]  = 1;
  ram[29580]  = 1;
  ram[29581]  = 1;
  ram[29582]  = 1;
  ram[29583]  = 1;
  ram[29584]  = 1;
  ram[29585]  = 1;
  ram[29586]  = 1;
  ram[29587]  = 1;
  ram[29588]  = 1;
  ram[29589]  = 1;
  ram[29590]  = 1;
  ram[29591]  = 1;
  ram[29592]  = 1;
  ram[29593]  = 1;
  ram[29594]  = 1;
  ram[29595]  = 1;
  ram[29596]  = 1;
  ram[29597]  = 1;
  ram[29598]  = 1;
  ram[29599]  = 1;
  ram[29600]  = 1;
  ram[29601]  = 1;
  ram[29602]  = 1;
  ram[29603]  = 1;
  ram[29604]  = 1;
  ram[29605]  = 1;
  ram[29606]  = 1;
  ram[29607]  = 1;
  ram[29608]  = 1;
  ram[29609]  = 1;
  ram[29610]  = 1;
  ram[29611]  = 1;
  ram[29612]  = 1;
  ram[29613]  = 1;
  ram[29614]  = 1;
  ram[29615]  = 1;
  ram[29616]  = 1;
  ram[29617]  = 1;
  ram[29618]  = 1;
  ram[29619]  = 1;
  ram[29620]  = 1;
  ram[29621]  = 1;
  ram[29622]  = 1;
  ram[29623]  = 1;
  ram[29624]  = 1;
  ram[29625]  = 1;
  ram[29626]  = 1;
  ram[29627]  = 1;
  ram[29628]  = 1;
  ram[29629]  = 1;
  ram[29630]  = 1;
  ram[29631]  = 1;
  ram[29632]  = 1;
  ram[29633]  = 1;
  ram[29634]  = 1;
  ram[29635]  = 1;
  ram[29636]  = 1;
  ram[29637]  = 1;
  ram[29638]  = 1;
  ram[29639]  = 1;
  ram[29640]  = 1;
  ram[29641]  = 1;
  ram[29642]  = 1;
  ram[29643]  = 1;
  ram[29644]  = 1;
  ram[29645]  = 1;
  ram[29646]  = 1;
  ram[29647]  = 1;
  ram[29648]  = 1;
  ram[29649]  = 1;
  ram[29650]  = 1;
  ram[29651]  = 1;
  ram[29652]  = 1;
  ram[29653]  = 1;
  ram[29654]  = 1;
  ram[29655]  = 1;
  ram[29656]  = 1;
  ram[29657]  = 1;
  ram[29658]  = 1;
  ram[29659]  = 1;
  ram[29660]  = 1;
  ram[29661]  = 1;
  ram[29662]  = 1;
  ram[29663]  = 1;
  ram[29664]  = 1;
  ram[29665]  = 1;
  ram[29666]  = 1;
  ram[29667]  = 1;
  ram[29668]  = 1;
  ram[29669]  = 1;
  ram[29670]  = 1;
  ram[29671]  = 1;
  ram[29672]  = 1;
  ram[29673]  = 1;
  ram[29674]  = 1;
  ram[29675]  = 1;
  ram[29676]  = 1;
  ram[29677]  = 1;
  ram[29678]  = 1;
  ram[29679]  = 1;
  ram[29680]  = 1;
  ram[29681]  = 1;
  ram[29682]  = 1;
  ram[29683]  = 1;
  ram[29684]  = 1;
  ram[29685]  = 1;
  ram[29686]  = 1;
  ram[29687]  = 1;
  ram[29688]  = 1;
  ram[29689]  = 1;
  ram[29690]  = 1;
  ram[29691]  = 1;
  ram[29692]  = 1;
  ram[29693]  = 1;
  ram[29694]  = 1;
  ram[29695]  = 1;
  ram[29696]  = 1;
  ram[29697]  = 1;
  ram[29698]  = 1;
  ram[29699]  = 1;
  ram[29700]  = 1;
  ram[29701]  = 1;
  ram[29702]  = 1;
  ram[29703]  = 1;
  ram[29704]  = 1;
  ram[29705]  = 1;
  ram[29706]  = 1;
  ram[29707]  = 1;
  ram[29708]  = 1;
  ram[29709]  = 1;
  ram[29710]  = 1;
  ram[29711]  = 1;
  ram[29712]  = 1;
  ram[29713]  = 1;
  ram[29714]  = 1;
  ram[29715]  = 1;
  ram[29716]  = 1;
  ram[29717]  = 1;
  ram[29718]  = 1;
  ram[29719]  = 1;
  ram[29720]  = 1;
  ram[29721]  = 1;
  ram[29722]  = 1;
  ram[29723]  = 1;
  ram[29724]  = 1;
  ram[29725]  = 1;
  ram[29726]  = 1;
  ram[29727]  = 1;
  ram[29728]  = 1;
  ram[29729]  = 1;
  ram[29730]  = 1;
  ram[29731]  = 1;
  ram[29732]  = 1;
  ram[29733]  = 1;
  ram[29734]  = 1;
  ram[29735]  = 1;
  ram[29736]  = 1;
  ram[29737]  = 1;
  ram[29738]  = 1;
  ram[29739]  = 1;
  ram[29740]  = 1;
  ram[29741]  = 1;
  ram[29742]  = 1;
  ram[29743]  = 1;
  ram[29744]  = 1;
  ram[29745]  = 1;
  ram[29746]  = 1;
  ram[29747]  = 1;
  ram[29748]  = 1;
  ram[29749]  = 1;
  ram[29750]  = 1;
  ram[29751]  = 1;
  ram[29752]  = 1;
  ram[29753]  = 1;
  ram[29754]  = 1;
  ram[29755]  = 1;
  ram[29756]  = 1;
  ram[29757]  = 1;
  ram[29758]  = 1;
  ram[29759]  = 1;
  ram[29760]  = 1;
  ram[29761]  = 1;
  ram[29762]  = 1;
  ram[29763]  = 1;
  ram[29764]  = 1;
  ram[29765]  = 1;
  ram[29766]  = 1;
  ram[29767]  = 1;
  ram[29768]  = 1;
  ram[29769]  = 1;
  ram[29770]  = 1;
  ram[29771]  = 1;
  ram[29772]  = 1;
  ram[29773]  = 1;
  ram[29774]  = 1;
  ram[29775]  = 1;
  ram[29776]  = 1;
  ram[29777]  = 1;
  ram[29778]  = 1;
  ram[29779]  = 1;
  ram[29780]  = 1;
  ram[29781]  = 1;
  ram[29782]  = 1;
  ram[29783]  = 1;
  ram[29784]  = 1;
  ram[29785]  = 1;
  ram[29786]  = 1;
  ram[29787]  = 1;
  ram[29788]  = 1;
  ram[29789]  = 1;
  ram[29790]  = 1;
  ram[29791]  = 1;
  ram[29792]  = 1;
  ram[29793]  = 1;
  ram[29794]  = 1;
  ram[29795]  = 1;
  ram[29796]  = 1;
  ram[29797]  = 1;
  ram[29798]  = 1;
  ram[29799]  = 1;
  ram[29800]  = 1;
  ram[29801]  = 1;
  ram[29802]  = 1;
  ram[29803]  = 1;
  ram[29804]  = 1;
  ram[29805]  = 1;
  ram[29806]  = 1;
  ram[29807]  = 1;
  ram[29808]  = 1;
  ram[29809]  = 1;
  ram[29810]  = 1;
  ram[29811]  = 1;
  ram[29812]  = 1;
  ram[29813]  = 1;
  ram[29814]  = 1;
  ram[29815]  = 1;
  ram[29816]  = 1;
  ram[29817]  = 1;
  ram[29818]  = 1;
  ram[29819]  = 1;
  ram[29820]  = 1;
  ram[29821]  = 1;
  ram[29822]  = 1;
  ram[29823]  = 1;
  ram[29824]  = 1;
  ram[29825]  = 1;
  ram[29826]  = 1;
  ram[29827]  = 1;
  ram[29828]  = 1;
  ram[29829]  = 1;
  ram[29830]  = 1;
  ram[29831]  = 1;
  ram[29832]  = 1;
  ram[29833]  = 1;
  ram[29834]  = 1;
  ram[29835]  = 1;
  ram[29836]  = 1;
  ram[29837]  = 1;
  ram[29838]  = 1;
  ram[29839]  = 1;
  ram[29840]  = 1;
  ram[29841]  = 1;
  ram[29842]  = 1;
  ram[29843]  = 1;
  ram[29844]  = 1;
  ram[29845]  = 1;
  ram[29846]  = 1;
  ram[29847]  = 1;
  ram[29848]  = 1;
  ram[29849]  = 1;
  ram[29850]  = 1;
  ram[29851]  = 1;
  ram[29852]  = 1;
  ram[29853]  = 1;
  ram[29854]  = 1;
  ram[29855]  = 1;
  ram[29856]  = 1;
  ram[29857]  = 1;
  ram[29858]  = 1;
  ram[29859]  = 1;
  ram[29860]  = 1;
  ram[29861]  = 1;
  ram[29862]  = 1;
  ram[29863]  = 1;
  ram[29864]  = 1;
  ram[29865]  = 1;
  ram[29866]  = 1;
  ram[29867]  = 1;
  ram[29868]  = 1;
  ram[29869]  = 1;
  ram[29870]  = 1;
  ram[29871]  = 1;
  ram[29872]  = 1;
  ram[29873]  = 1;
  ram[29874]  = 1;
  ram[29875]  = 1;
  ram[29876]  = 1;
  ram[29877]  = 1;
  ram[29878]  = 1;
  ram[29879]  = 1;
  ram[29880]  = 1;
  ram[29881]  = 1;
  ram[29882]  = 1;
  ram[29883]  = 1;
  ram[29884]  = 1;
  ram[29885]  = 1;
  ram[29886]  = 1;
  ram[29887]  = 1;
  ram[29888]  = 1;
  ram[29889]  = 1;
  ram[29890]  = 1;
  ram[29891]  = 1;
  ram[29892]  = 1;
  ram[29893]  = 1;
  ram[29894]  = 1;
  ram[29895]  = 1;
  ram[29896]  = 1;
  ram[29897]  = 1;
  ram[29898]  = 1;
  ram[29899]  = 1;
  ram[29900]  = 1;
  ram[29901]  = 1;
  ram[29902]  = 1;
  ram[29903]  = 1;
  ram[29904]  = 1;
  ram[29905]  = 1;
  ram[29906]  = 1;
  ram[29907]  = 1;
  ram[29908]  = 1;
  ram[29909]  = 1;
  ram[29910]  = 1;
  ram[29911]  = 1;
  ram[29912]  = 1;
  ram[29913]  = 1;
  ram[29914]  = 1;
  ram[29915]  = 1;
  ram[29916]  = 1;
  ram[29917]  = 1;
  ram[29918]  = 1;
  ram[29919]  = 1;
  ram[29920]  = 1;
  ram[29921]  = 1;
  ram[29922]  = 1;
  ram[29923]  = 1;
  ram[29924]  = 1;
  ram[29925]  = 1;
  ram[29926]  = 1;
  ram[29927]  = 1;
  ram[29928]  = 1;
  ram[29929]  = 1;
  ram[29930]  = 1;
  ram[29931]  = 1;
  ram[29932]  = 1;
  ram[29933]  = 1;
  ram[29934]  = 1;
  ram[29935]  = 1;
  ram[29936]  = 1;
  ram[29937]  = 1;
  ram[29938]  = 1;
  ram[29939]  = 1;
  ram[29940]  = 1;
  ram[29941]  = 1;
  ram[29942]  = 1;
  ram[29943]  = 1;
  ram[29944]  = 1;
  ram[29945]  = 1;
  ram[29946]  = 1;
  ram[29947]  = 1;
  ram[29948]  = 1;
  ram[29949]  = 1;
  ram[29950]  = 1;
  ram[29951]  = 1;
  ram[29952]  = 1;
  ram[29953]  = 1;
  ram[29954]  = 1;
  ram[29955]  = 1;
  ram[29956]  = 1;
  ram[29957]  = 1;
  ram[29958]  = 1;
  ram[29959]  = 1;
  ram[29960]  = 1;
  ram[29961]  = 1;
  ram[29962]  = 1;
  ram[29963]  = 1;
  ram[29964]  = 1;
  ram[29965]  = 1;
  ram[29966]  = 1;
  ram[29967]  = 1;
  ram[29968]  = 1;
  ram[29969]  = 1;
  ram[29970]  = 1;
  ram[29971]  = 1;
  ram[29972]  = 1;
  ram[29973]  = 1;
  ram[29974]  = 1;
  ram[29975]  = 1;
  ram[29976]  = 1;
  ram[29977]  = 1;
  ram[29978]  = 1;
  ram[29979]  = 1;
  ram[29980]  = 1;
  ram[29981]  = 1;
  ram[29982]  = 1;
  ram[29983]  = 1;
  ram[29984]  = 1;
  ram[29985]  = 1;
  ram[29986]  = 1;
  ram[29987]  = 1;
  ram[29988]  = 1;
  ram[29989]  = 1;
  ram[29990]  = 1;
  ram[29991]  = 1;
  ram[29992]  = 1;
  ram[29993]  = 1;
  ram[29994]  = 1;
  ram[29995]  = 1;
  ram[29996]  = 1;
  ram[29997]  = 1;
  ram[29998]  = 1;
  ram[29999]  = 1;
  ram[30000]  = 1;
  ram[30001]  = 1;
  ram[30002]  = 1;
  ram[30003]  = 1;
  ram[30004]  = 1;
  ram[30005]  = 1;
  ram[30006]  = 1;
  ram[30007]  = 1;
  ram[30008]  = 1;
  ram[30009]  = 1;
  ram[30010]  = 1;
  ram[30011]  = 1;
  ram[30012]  = 1;
  ram[30013]  = 1;
  ram[30014]  = 1;
  ram[30015]  = 1;
  ram[30016]  = 1;
  ram[30017]  = 1;
  ram[30018]  = 1;
  ram[30019]  = 1;
  ram[30020]  = 1;
  ram[30021]  = 1;
  ram[30022]  = 1;
  ram[30023]  = 1;
  ram[30024]  = 1;
  ram[30025]  = 1;
  ram[30026]  = 1;
  ram[30027]  = 1;
  ram[30028]  = 1;
  ram[30029]  = 1;
  ram[30030]  = 1;
  ram[30031]  = 1;
  ram[30032]  = 1;
  ram[30033]  = 1;
  ram[30034]  = 1;
  ram[30035]  = 1;
  ram[30036]  = 1;
  ram[30037]  = 1;
  ram[30038]  = 1;
  ram[30039]  = 1;
  ram[30040]  = 1;
  ram[30041]  = 1;
  ram[30042]  = 1;
  ram[30043]  = 1;
  ram[30044]  = 1;
  ram[30045]  = 1;
  ram[30046]  = 1;
  ram[30047]  = 1;
  ram[30048]  = 1;
  ram[30049]  = 1;
  ram[30050]  = 1;
  ram[30051]  = 1;
  ram[30052]  = 1;
  ram[30053]  = 1;
  ram[30054]  = 1;
  ram[30055]  = 1;
  ram[30056]  = 1;
  ram[30057]  = 1;
  ram[30058]  = 1;
  ram[30059]  = 1;
  ram[30060]  = 1;
  ram[30061]  = 1;
  ram[30062]  = 1;
  ram[30063]  = 1;
  ram[30064]  = 1;
  ram[30065]  = 1;
  ram[30066]  = 1;
  ram[30067]  = 1;
  ram[30068]  = 1;
  ram[30069]  = 1;
  ram[30070]  = 1;
  ram[30071]  = 1;
  ram[30072]  = 1;
  ram[30073]  = 1;
  ram[30074]  = 1;
  ram[30075]  = 1;
  ram[30076]  = 1;
  ram[30077]  = 1;
  ram[30078]  = 1;
  ram[30079]  = 1;
  ram[30080]  = 1;
  ram[30081]  = 1;
  ram[30082]  = 1;
  ram[30083]  = 1;
  ram[30084]  = 1;
  ram[30085]  = 1;
  ram[30086]  = 1;
  ram[30087]  = 1;
  ram[30088]  = 1;
  ram[30089]  = 1;
  ram[30090]  = 1;
  ram[30091]  = 1;
  ram[30092]  = 1;
  ram[30093]  = 1;
  ram[30094]  = 1;
  ram[30095]  = 1;
  ram[30096]  = 1;
  ram[30097]  = 1;
  ram[30098]  = 1;
  ram[30099]  = 1;
  ram[30100]  = 1;
  ram[30101]  = 1;
  ram[30102]  = 1;
  ram[30103]  = 1;
  ram[30104]  = 1;
  ram[30105]  = 1;
  ram[30106]  = 1;
  ram[30107]  = 1;
  ram[30108]  = 1;
  ram[30109]  = 1;
  ram[30110]  = 1;
  ram[30111]  = 1;
  ram[30112]  = 1;
  ram[30113]  = 1;
  ram[30114]  = 1;
  ram[30115]  = 1;
  ram[30116]  = 1;
  ram[30117]  = 1;
  ram[30118]  = 1;
  ram[30119]  = 1;
  ram[30120]  = 1;
  ram[30121]  = 1;
  ram[30122]  = 1;
  ram[30123]  = 1;
  ram[30124]  = 1;
  ram[30125]  = 1;
  ram[30126]  = 1;
  ram[30127]  = 1;
  ram[30128]  = 1;
  ram[30129]  = 1;
  ram[30130]  = 1;
  ram[30131]  = 1;
  ram[30132]  = 1;
  ram[30133]  = 1;
  ram[30134]  = 1;
  ram[30135]  = 1;
  ram[30136]  = 1;
  ram[30137]  = 1;
  ram[30138]  = 1;
  ram[30139]  = 1;
  ram[30140]  = 1;
  ram[30141]  = 1;
  ram[30142]  = 1;
  ram[30143]  = 1;
  ram[30144]  = 1;
  ram[30145]  = 1;
  ram[30146]  = 1;
  ram[30147]  = 1;
  ram[30148]  = 1;
  ram[30149]  = 1;
  ram[30150]  = 1;
  ram[30151]  = 1;
  ram[30152]  = 1;
  ram[30153]  = 1;
  ram[30154]  = 1;
  ram[30155]  = 1;
  ram[30156]  = 1;
  ram[30157]  = 1;
  ram[30158]  = 1;
  ram[30159]  = 1;
  ram[30160]  = 1;
  ram[30161]  = 1;
  ram[30162]  = 1;
  ram[30163]  = 1;
  ram[30164]  = 1;
  ram[30165]  = 1;
  ram[30166]  = 1;
  ram[30167]  = 1;
  ram[30168]  = 1;
  ram[30169]  = 1;
  ram[30170]  = 1;
  ram[30171]  = 1;
  ram[30172]  = 1;
  ram[30173]  = 1;
  ram[30174]  = 1;
  ram[30175]  = 1;
  ram[30176]  = 1;
  ram[30177]  = 1;
  ram[30178]  = 1;
  ram[30179]  = 1;
  ram[30180]  = 1;
  ram[30181]  = 1;
  ram[30182]  = 1;
  ram[30183]  = 1;
  ram[30184]  = 1;
  ram[30185]  = 1;
  ram[30186]  = 1;
  ram[30187]  = 1;
  ram[30188]  = 1;
  ram[30189]  = 1;
  ram[30190]  = 1;
  ram[30191]  = 1;
  ram[30192]  = 1;
  ram[30193]  = 1;
  ram[30194]  = 1;
  ram[30195]  = 1;
  ram[30196]  = 1;
  ram[30197]  = 1;
  ram[30198]  = 1;
  ram[30199]  = 1;
  ram[30200]  = 1;
  ram[30201]  = 1;
  ram[30202]  = 1;
  ram[30203]  = 1;
  ram[30204]  = 1;
  ram[30205]  = 1;
  ram[30206]  = 1;
  ram[30207]  = 1;
  ram[30208]  = 1;
  ram[30209]  = 1;
  ram[30210]  = 1;
  ram[30211]  = 1;
  ram[30212]  = 1;
  ram[30213]  = 1;
  ram[30214]  = 1;
  ram[30215]  = 1;
  ram[30216]  = 1;
  ram[30217]  = 1;
  ram[30218]  = 1;
  ram[30219]  = 1;
  ram[30220]  = 1;
  ram[30221]  = 1;
  ram[30222]  = 1;
  ram[30223]  = 1;
  ram[30224]  = 1;
  ram[30225]  = 1;
  ram[30226]  = 1;
  ram[30227]  = 1;
  ram[30228]  = 1;
  ram[30229]  = 1;
  ram[30230]  = 1;
  ram[30231]  = 1;
  ram[30232]  = 1;
  ram[30233]  = 1;
  ram[30234]  = 1;
  ram[30235]  = 1;
  ram[30236]  = 1;
  ram[30237]  = 1;
  ram[30238]  = 1;
  ram[30239]  = 1;
  ram[30240]  = 1;
  ram[30241]  = 1;
  ram[30242]  = 1;
  ram[30243]  = 1;
  ram[30244]  = 1;
  ram[30245]  = 1;
  ram[30246]  = 1;
  ram[30247]  = 1;
  ram[30248]  = 1;
  ram[30249]  = 1;
  ram[30250]  = 1;
  ram[30251]  = 1;
  ram[30252]  = 1;
  ram[30253]  = 1;
  ram[30254]  = 1;
  ram[30255]  = 1;
  ram[30256]  = 1;
  ram[30257]  = 1;
  ram[30258]  = 1;
  ram[30259]  = 1;
  ram[30260]  = 1;
  ram[30261]  = 1;
  ram[30262]  = 1;
  ram[30263]  = 1;
  ram[30264]  = 1;
  ram[30265]  = 1;
  ram[30266]  = 1;
  ram[30267]  = 1;
  ram[30268]  = 1;
  ram[30269]  = 1;
  ram[30270]  = 1;
  ram[30271]  = 1;
  ram[30272]  = 1;
  ram[30273]  = 1;
  ram[30274]  = 1;
  ram[30275]  = 1;
  ram[30276]  = 1;
  ram[30277]  = 1;
  ram[30278]  = 1;
  ram[30279]  = 1;
  ram[30280]  = 1;
  ram[30281]  = 1;
  ram[30282]  = 1;
  ram[30283]  = 1;
  ram[30284]  = 1;
  ram[30285]  = 1;
  ram[30286]  = 1;
  ram[30287]  = 1;
  ram[30288]  = 1;
  ram[30289]  = 1;
  ram[30290]  = 1;
  ram[30291]  = 1;
  ram[30292]  = 1;
  ram[30293]  = 1;
  ram[30294]  = 1;
  ram[30295]  = 1;
  ram[30296]  = 1;
  ram[30297]  = 1;
  ram[30298]  = 1;
  ram[30299]  = 1;
  ram[30300]  = 1;
  ram[30301]  = 1;
  ram[30302]  = 1;
  ram[30303]  = 1;
  ram[30304]  = 1;
  ram[30305]  = 1;
  ram[30306]  = 1;
  ram[30307]  = 1;
  ram[30308]  = 1;
  ram[30309]  = 1;
  ram[30310]  = 1;
  ram[30311]  = 1;
  ram[30312]  = 1;
  ram[30313]  = 1;
  ram[30314]  = 1;
  ram[30315]  = 1;
  ram[30316]  = 1;
  ram[30317]  = 1;
  ram[30318]  = 1;
  ram[30319]  = 1;
  ram[30320]  = 1;
  ram[30321]  = 1;
  ram[30322]  = 1;
  ram[30323]  = 1;
  ram[30324]  = 1;
  ram[30325]  = 1;
  ram[30326]  = 1;
  ram[30327]  = 1;
  ram[30328]  = 1;
  ram[30329]  = 1;
  ram[30330]  = 1;
  ram[30331]  = 1;
  ram[30332]  = 1;
  ram[30333]  = 1;
  ram[30334]  = 1;
  ram[30335]  = 1;
  ram[30336]  = 1;
  ram[30337]  = 1;
  ram[30338]  = 1;
  ram[30339]  = 1;
  ram[30340]  = 1;
  ram[30341]  = 1;
  ram[30342]  = 1;
  ram[30343]  = 1;
  ram[30344]  = 1;
  ram[30345]  = 1;
  ram[30346]  = 1;
  ram[30347]  = 1;
  ram[30348]  = 1;
  ram[30349]  = 1;
  ram[30350]  = 1;
  ram[30351]  = 1;
  ram[30352]  = 1;
  ram[30353]  = 1;
  ram[30354]  = 1;
  ram[30355]  = 1;
  ram[30356]  = 1;
  ram[30357]  = 1;
  ram[30358]  = 1;
  ram[30359]  = 1;
  ram[30360]  = 1;
  ram[30361]  = 1;
  ram[30362]  = 1;
  ram[30363]  = 1;
  ram[30364]  = 1;
  ram[30365]  = 1;
  ram[30366]  = 1;
  ram[30367]  = 1;
  ram[30368]  = 1;
  ram[30369]  = 1;
  ram[30370]  = 1;
  ram[30371]  = 1;
  ram[30372]  = 1;
  ram[30373]  = 1;
  ram[30374]  = 1;
  ram[30375]  = 1;
  ram[30376]  = 1;
  ram[30377]  = 1;
  ram[30378]  = 1;
  ram[30379]  = 1;
  ram[30380]  = 1;
  ram[30381]  = 1;
  ram[30382]  = 1;
  ram[30383]  = 1;
  ram[30384]  = 1;
  ram[30385]  = 1;
  ram[30386]  = 1;
  ram[30387]  = 1;
  ram[30388]  = 1;
  ram[30389]  = 1;
  ram[30390]  = 1;
  ram[30391]  = 1;
  ram[30392]  = 1;
  ram[30393]  = 1;
  ram[30394]  = 1;
  ram[30395]  = 1;
  ram[30396]  = 1;
  ram[30397]  = 1;
  ram[30398]  = 1;
  ram[30399]  = 1;
  ram[30400]  = 1;
  ram[30401]  = 1;
  ram[30402]  = 1;
  ram[30403]  = 1;
  ram[30404]  = 1;
  ram[30405]  = 1;
  ram[30406]  = 1;
  ram[30407]  = 1;
  ram[30408]  = 1;
  ram[30409]  = 1;
  ram[30410]  = 1;
  ram[30411]  = 1;
  ram[30412]  = 1;
  ram[30413]  = 1;
  ram[30414]  = 1;
  ram[30415]  = 1;
  ram[30416]  = 1;
  ram[30417]  = 1;
  ram[30418]  = 1;
  ram[30419]  = 1;
  ram[30420]  = 1;
  ram[30421]  = 1;
  ram[30422]  = 1;
  ram[30423]  = 1;
  ram[30424]  = 1;
  ram[30425]  = 1;
  ram[30426]  = 1;
  ram[30427]  = 1;
  ram[30428]  = 1;
  ram[30429]  = 1;
  ram[30430]  = 1;
  ram[30431]  = 1;
  ram[30432]  = 1;
  ram[30433]  = 1;
  ram[30434]  = 1;
  ram[30435]  = 1;
  ram[30436]  = 1;
  ram[30437]  = 1;
  ram[30438]  = 1;
  ram[30439]  = 1;
  ram[30440]  = 1;
  ram[30441]  = 1;
  ram[30442]  = 1;
  ram[30443]  = 1;
  ram[30444]  = 1;
  ram[30445]  = 1;
  ram[30446]  = 1;
  ram[30447]  = 1;
  ram[30448]  = 1;
  ram[30449]  = 1;
  ram[30450]  = 1;
  ram[30451]  = 1;
  ram[30452]  = 1;
  ram[30453]  = 1;
  ram[30454]  = 1;
  ram[30455]  = 1;
  ram[30456]  = 1;
  ram[30457]  = 1;
  ram[30458]  = 1;
  ram[30459]  = 1;
  ram[30460]  = 1;
  ram[30461]  = 1;
  ram[30462]  = 1;
  ram[30463]  = 1;
  ram[30464]  = 1;
  ram[30465]  = 1;
  ram[30466]  = 1;
  ram[30467]  = 1;
  ram[30468]  = 1;
  ram[30469]  = 1;
  ram[30470]  = 1;
  ram[30471]  = 1;
  ram[30472]  = 1;
  ram[30473]  = 1;
  ram[30474]  = 1;
  ram[30475]  = 1;
  ram[30476]  = 1;
  ram[30477]  = 1;
  ram[30478]  = 1;
  ram[30479]  = 1;
  ram[30480]  = 1;
  ram[30481]  = 1;
  ram[30482]  = 1;
  ram[30483]  = 1;
  ram[30484]  = 1;
  ram[30485]  = 1;
  ram[30486]  = 1;
  ram[30487]  = 1;
  ram[30488]  = 1;
  ram[30489]  = 1;
  ram[30490]  = 1;
  ram[30491]  = 1;
  ram[30492]  = 1;
  ram[30493]  = 1;
  ram[30494]  = 1;
  ram[30495]  = 1;
  ram[30496]  = 1;
  ram[30497]  = 1;
  ram[30498]  = 1;
  ram[30499]  = 1;
  ram[30500]  = 1;
  ram[30501]  = 1;
  ram[30502]  = 1;
  ram[30503]  = 1;
  ram[30504]  = 1;
  ram[30505]  = 1;
  ram[30506]  = 1;
  ram[30507]  = 1;
  ram[30508]  = 1;
  ram[30509]  = 1;
  ram[30510]  = 1;
  ram[30511]  = 1;
  ram[30512]  = 1;
  ram[30513]  = 1;
  ram[30514]  = 1;
  ram[30515]  = 1;
  ram[30516]  = 1;
  ram[30517]  = 1;
  ram[30518]  = 1;
  ram[30519]  = 1;
  ram[30520]  = 1;
  ram[30521]  = 1;
  ram[30522]  = 1;
  ram[30523]  = 1;
  ram[30524]  = 1;
  ram[30525]  = 1;
  ram[30526]  = 1;
  ram[30527]  = 1;
  ram[30528]  = 1;
  ram[30529]  = 1;
  ram[30530]  = 1;
  ram[30531]  = 1;
  ram[30532]  = 1;
  ram[30533]  = 1;
  ram[30534]  = 1;
  ram[30535]  = 1;
  ram[30536]  = 1;
  ram[30537]  = 1;
  ram[30538]  = 1;
  ram[30539]  = 1;
  ram[30540]  = 1;
  ram[30541]  = 1;
  ram[30542]  = 1;
  ram[30543]  = 1;
  ram[30544]  = 1;
  ram[30545]  = 1;
  ram[30546]  = 1;
  ram[30547]  = 1;
  ram[30548]  = 1;
  ram[30549]  = 1;
  ram[30550]  = 1;
  ram[30551]  = 1;
  ram[30552]  = 1;
  ram[30553]  = 1;
  ram[30554]  = 1;
  ram[30555]  = 1;
  ram[30556]  = 1;
  ram[30557]  = 1;
  ram[30558]  = 1;
  ram[30559]  = 1;
  ram[30560]  = 1;
  ram[30561]  = 1;
  ram[30562]  = 1;
  ram[30563]  = 1;
  ram[30564]  = 1;
  ram[30565]  = 1;
  ram[30566]  = 1;
  ram[30567]  = 1;
  ram[30568]  = 1;
  ram[30569]  = 1;
  ram[30570]  = 1;
  ram[30571]  = 1;
  ram[30572]  = 1;
  ram[30573]  = 1;
  ram[30574]  = 1;
  ram[30575]  = 1;
  ram[30576]  = 1;
  ram[30577]  = 1;
  ram[30578]  = 1;
  ram[30579]  = 1;
  ram[30580]  = 1;
  ram[30581]  = 1;
  ram[30582]  = 1;
  ram[30583]  = 1;
  ram[30584]  = 1;
  ram[30585]  = 1;
  ram[30586]  = 1;
  ram[30587]  = 1;
  ram[30588]  = 1;
  ram[30589]  = 1;
  ram[30590]  = 1;
  ram[30591]  = 1;
  ram[30592]  = 1;
  ram[30593]  = 1;
  ram[30594]  = 1;
  ram[30595]  = 1;
  ram[30596]  = 1;
  ram[30597]  = 1;
  ram[30598]  = 1;
  ram[30599]  = 1;
  ram[30600]  = 1;
  ram[30601]  = 1;
  ram[30602]  = 1;
  ram[30603]  = 1;
  ram[30604]  = 1;
  ram[30605]  = 1;
  ram[30606]  = 1;
  ram[30607]  = 1;
  ram[30608]  = 1;
  ram[30609]  = 1;
  ram[30610]  = 1;
  ram[30611]  = 1;
  ram[30612]  = 1;
  ram[30613]  = 1;
  ram[30614]  = 1;
  ram[30615]  = 1;
  ram[30616]  = 1;
  ram[30617]  = 1;
  ram[30618]  = 1;
  ram[30619]  = 1;
  ram[30620]  = 1;
  ram[30621]  = 1;
  ram[30622]  = 1;
  ram[30623]  = 1;
  ram[30624]  = 1;
  ram[30625]  = 1;
  ram[30626]  = 1;
  ram[30627]  = 1;
  ram[30628]  = 1;
  ram[30629]  = 1;
  ram[30630]  = 1;
  ram[30631]  = 1;
  ram[30632]  = 1;
  ram[30633]  = 1;
  ram[30634]  = 1;
  ram[30635]  = 1;
  ram[30636]  = 1;
  ram[30637]  = 1;
  ram[30638]  = 1;
  ram[30639]  = 1;
  ram[30640]  = 1;
  ram[30641]  = 1;
  ram[30642]  = 1;
  ram[30643]  = 1;
  ram[30644]  = 1;
  ram[30645]  = 1;
  ram[30646]  = 1;
  ram[30647]  = 1;
  ram[30648]  = 1;
  ram[30649]  = 1;
  ram[30650]  = 1;
  ram[30651]  = 1;
  ram[30652]  = 1;
  ram[30653]  = 1;
  ram[30654]  = 1;
  ram[30655]  = 1;
  ram[30656]  = 1;
  ram[30657]  = 1;
  ram[30658]  = 1;
  ram[30659]  = 1;
  ram[30660]  = 1;
  ram[30661]  = 1;
  ram[30662]  = 1;
  ram[30663]  = 1;
  ram[30664]  = 1;
  ram[30665]  = 1;
  ram[30666]  = 1;
  ram[30667]  = 1;
  ram[30668]  = 1;
  ram[30669]  = 1;
  ram[30670]  = 1;
  ram[30671]  = 1;
  ram[30672]  = 1;
  ram[30673]  = 1;
  ram[30674]  = 1;
  ram[30675]  = 1;
  ram[30676]  = 1;
  ram[30677]  = 1;
  ram[30678]  = 1;
  ram[30679]  = 1;
  ram[30680]  = 1;
  ram[30681]  = 1;
  ram[30682]  = 1;
  ram[30683]  = 1;
  ram[30684]  = 1;
  ram[30685]  = 1;
  ram[30686]  = 1;
  ram[30687]  = 1;
  ram[30688]  = 1;
  ram[30689]  = 1;
  ram[30690]  = 1;
  ram[30691]  = 1;
  ram[30692]  = 1;
  ram[30693]  = 1;
  ram[30694]  = 1;
  ram[30695]  = 1;
  ram[30696]  = 1;
  ram[30697]  = 1;
  ram[30698]  = 1;
  ram[30699]  = 1;
  ram[30700]  = 1;
  ram[30701]  = 1;
  ram[30702]  = 1;
  ram[30703]  = 1;
  ram[30704]  = 1;
  ram[30705]  = 1;
  ram[30706]  = 1;
  ram[30707]  = 1;
  ram[30708]  = 1;
  ram[30709]  = 1;
  ram[30710]  = 1;
  ram[30711]  = 1;
  ram[30712]  = 1;
  ram[30713]  = 1;
  ram[30714]  = 1;
  ram[30715]  = 1;
  ram[30716]  = 1;
  ram[30717]  = 1;
  ram[30718]  = 1;
  ram[30719]  = 1;
  ram[30720]  = 1;
  ram[30721]  = 1;
  ram[30722]  = 1;
  ram[30723]  = 1;
  ram[30724]  = 1;
  ram[30725]  = 1;
  ram[30726]  = 1;
  ram[30727]  = 1;
  ram[30728]  = 1;
  ram[30729]  = 1;
  ram[30730]  = 1;
  ram[30731]  = 1;
  ram[30732]  = 1;
  ram[30733]  = 1;
  ram[30734]  = 1;
  ram[30735]  = 1;
  ram[30736]  = 1;
  ram[30737]  = 1;
  ram[30738]  = 1;
  ram[30739]  = 1;
  ram[30740]  = 1;
  ram[30741]  = 1;
  ram[30742]  = 1;
  ram[30743]  = 1;
  ram[30744]  = 1;
  ram[30745]  = 1;
  ram[30746]  = 1;
  ram[30747]  = 1;
  ram[30748]  = 1;
  ram[30749]  = 1;
  ram[30750]  = 1;
  ram[30751]  = 1;
  ram[30752]  = 1;
  ram[30753]  = 1;
  ram[30754]  = 1;
  ram[30755]  = 1;
  ram[30756]  = 1;
  ram[30757]  = 1;
  ram[30758]  = 1;
  ram[30759]  = 1;
  ram[30760]  = 1;
  ram[30761]  = 1;
  ram[30762]  = 1;
  ram[30763]  = 1;
  ram[30764]  = 1;
  ram[30765]  = 1;
  ram[30766]  = 1;
  ram[30767]  = 1;
  ram[30768]  = 1;
  ram[30769]  = 1;
  ram[30770]  = 1;
  ram[30771]  = 1;
  ram[30772]  = 1;
  ram[30773]  = 1;
  ram[30774]  = 1;
  ram[30775]  = 1;
  ram[30776]  = 1;
  ram[30777]  = 1;
  ram[30778]  = 1;
  ram[30779]  = 1;
  ram[30780]  = 1;
  ram[30781]  = 1;
  ram[30782]  = 1;
  ram[30783]  = 1;
  ram[30784]  = 1;
  ram[30785]  = 1;
  ram[30786]  = 1;
  ram[30787]  = 1;
  ram[30788]  = 1;
  ram[30789]  = 1;
  ram[30790]  = 1;
  ram[30791]  = 1;
  ram[30792]  = 1;
  ram[30793]  = 1;
  ram[30794]  = 1;
  ram[30795]  = 1;
  ram[30796]  = 1;
  ram[30797]  = 1;
  ram[30798]  = 1;
  ram[30799]  = 1;
  ram[30800]  = 1;
  ram[30801]  = 1;
  ram[30802]  = 1;
  ram[30803]  = 1;
  ram[30804]  = 1;
  ram[30805]  = 1;
  ram[30806]  = 1;
  ram[30807]  = 1;
  ram[30808]  = 1;
  ram[30809]  = 1;
  ram[30810]  = 1;
  ram[30811]  = 1;
  ram[30812]  = 1;
  ram[30813]  = 1;
  ram[30814]  = 1;
  ram[30815]  = 1;
  ram[30816]  = 1;
  ram[30817]  = 1;
  ram[30818]  = 1;
  ram[30819]  = 1;
  ram[30820]  = 1;
  ram[30821]  = 1;
  ram[30822]  = 1;
  ram[30823]  = 1;
  ram[30824]  = 1;
  ram[30825]  = 1;
  ram[30826]  = 1;
  ram[30827]  = 1;
  ram[30828]  = 1;
  ram[30829]  = 1;
  ram[30830]  = 1;
  ram[30831]  = 1;
  ram[30832]  = 1;
  ram[30833]  = 1;
  ram[30834]  = 1;
  ram[30835]  = 1;
  ram[30836]  = 1;
  ram[30837]  = 1;
  ram[30838]  = 1;
  ram[30839]  = 1;
  ram[30840]  = 1;
  ram[30841]  = 1;
  ram[30842]  = 1;
  ram[30843]  = 1;
  ram[30844]  = 1;
  ram[30845]  = 1;
  ram[30846]  = 1;
  ram[30847]  = 1;
  ram[30848]  = 1;
  ram[30849]  = 1;
  ram[30850]  = 1;
  ram[30851]  = 1;
  ram[30852]  = 1;
  ram[30853]  = 1;
  ram[30854]  = 1;
  ram[30855]  = 1;
  ram[30856]  = 1;
  ram[30857]  = 1;
  ram[30858]  = 1;
  ram[30859]  = 1;
  ram[30860]  = 1;
  ram[30861]  = 1;
  ram[30862]  = 1;
  ram[30863]  = 1;
  ram[30864]  = 1;
  ram[30865]  = 1;
  ram[30866]  = 1;
  ram[30867]  = 1;
  ram[30868]  = 1;
  ram[30869]  = 1;
  ram[30870]  = 1;
  ram[30871]  = 1;
  ram[30872]  = 1;
  ram[30873]  = 1;
  ram[30874]  = 1;
  ram[30875]  = 1;
  ram[30876]  = 1;
  ram[30877]  = 1;
  ram[30878]  = 1;
  ram[30879]  = 1;
  ram[30880]  = 1;
  ram[30881]  = 1;
  ram[30882]  = 1;
  ram[30883]  = 1;
  ram[30884]  = 1;
  ram[30885]  = 1;
  ram[30886]  = 1;
  ram[30887]  = 1;
  ram[30888]  = 1;
  ram[30889]  = 1;
  ram[30890]  = 1;
  ram[30891]  = 1;
  ram[30892]  = 1;
  ram[30893]  = 1;
  ram[30894]  = 1;
  ram[30895]  = 1;
  ram[30896]  = 1;
  ram[30897]  = 1;
  ram[30898]  = 1;
  ram[30899]  = 1;
  ram[30900]  = 1;
  ram[30901]  = 1;
  ram[30902]  = 1;
  ram[30903]  = 1;
  ram[30904]  = 1;
  ram[30905]  = 1;
  ram[30906]  = 1;
  ram[30907]  = 1;
  ram[30908]  = 1;
  ram[30909]  = 1;
  ram[30910]  = 1;
  ram[30911]  = 1;
  ram[30912]  = 1;
  ram[30913]  = 1;
  ram[30914]  = 1;
  ram[30915]  = 1;
  ram[30916]  = 1;
  ram[30917]  = 1;
  ram[30918]  = 1;
  ram[30919]  = 1;
  ram[30920]  = 1;
  ram[30921]  = 1;
  ram[30922]  = 1;
  ram[30923]  = 1;
  ram[30924]  = 1;
  ram[30925]  = 1;
  ram[30926]  = 1;
  ram[30927]  = 1;
  ram[30928]  = 1;
  ram[30929]  = 1;
  ram[30930]  = 1;
  ram[30931]  = 1;
  ram[30932]  = 1;
  ram[30933]  = 1;
  ram[30934]  = 1;
  ram[30935]  = 1;
  ram[30936]  = 1;
  ram[30937]  = 1;
  ram[30938]  = 1;
  ram[30939]  = 1;
  ram[30940]  = 1;
  ram[30941]  = 1;
  ram[30942]  = 1;
  ram[30943]  = 1;
  ram[30944]  = 1;
  ram[30945]  = 1;
  ram[30946]  = 1;
  ram[30947]  = 1;
  ram[30948]  = 1;
  ram[30949]  = 1;
  ram[30950]  = 1;
  ram[30951]  = 1;
  ram[30952]  = 1;
  ram[30953]  = 1;
  ram[30954]  = 1;
  ram[30955]  = 1;
  ram[30956]  = 1;
  ram[30957]  = 1;
  ram[30958]  = 1;
  ram[30959]  = 1;
  ram[30960]  = 1;
  ram[30961]  = 1;
  ram[30962]  = 1;
  ram[30963]  = 1;
  ram[30964]  = 1;
  ram[30965]  = 1;
  ram[30966]  = 1;
  ram[30967]  = 1;
  ram[30968]  = 1;
  ram[30969]  = 1;
  ram[30970]  = 1;
  ram[30971]  = 1;
  ram[30972]  = 1;
  ram[30973]  = 1;
  ram[30974]  = 1;
  ram[30975]  = 1;
  ram[30976]  = 1;
  ram[30977]  = 1;
  ram[30978]  = 1;
  ram[30979]  = 1;
  ram[30980]  = 1;
  ram[30981]  = 1;
  ram[30982]  = 1;
  ram[30983]  = 1;
  ram[30984]  = 1;
  ram[30985]  = 1;
  ram[30986]  = 1;
  ram[30987]  = 1;
  ram[30988]  = 1;
  ram[30989]  = 1;
  ram[30990]  = 1;
  ram[30991]  = 1;
  ram[30992]  = 1;
  ram[30993]  = 1;
  ram[30994]  = 1;
  ram[30995]  = 1;
  ram[30996]  = 1;
  ram[30997]  = 1;
  ram[30998]  = 1;
  ram[30999]  = 1;
  ram[31000]  = 1;
  ram[31001]  = 1;
  ram[31002]  = 1;
  ram[31003]  = 1;
  ram[31004]  = 1;
  ram[31005]  = 1;
  ram[31006]  = 1;
  ram[31007]  = 1;
  ram[31008]  = 1;
  ram[31009]  = 1;
  ram[31010]  = 1;
  ram[31011]  = 1;
  ram[31012]  = 1;
  ram[31013]  = 1;
  ram[31014]  = 1;
  ram[31015]  = 1;
  ram[31016]  = 1;
  ram[31017]  = 1;
  ram[31018]  = 1;
  ram[31019]  = 1;
  ram[31020]  = 1;
  ram[31021]  = 1;
  ram[31022]  = 1;
  ram[31023]  = 1;
  ram[31024]  = 1;
  ram[31025]  = 1;
  ram[31026]  = 1;
  ram[31027]  = 1;
  ram[31028]  = 1;
  ram[31029]  = 1;
  ram[31030]  = 1;
  ram[31031]  = 1;
  ram[31032]  = 1;
  ram[31033]  = 1;
  ram[31034]  = 1;
  ram[31035]  = 1;
  ram[31036]  = 1;
  ram[31037]  = 1;
  ram[31038]  = 1;
  ram[31039]  = 1;
  ram[31040]  = 1;
  ram[31041]  = 1;
  ram[31042]  = 1;
  ram[31043]  = 1;
  ram[31044]  = 1;
  ram[31045]  = 1;
  ram[31046]  = 1;
  ram[31047]  = 1;
  ram[31048]  = 1;
  ram[31049]  = 1;
  ram[31050]  = 1;
  ram[31051]  = 1;
  ram[31052]  = 1;
  ram[31053]  = 1;
  ram[31054]  = 1;
  ram[31055]  = 1;
  ram[31056]  = 1;
  ram[31057]  = 1;
  ram[31058]  = 1;
  ram[31059]  = 1;
  ram[31060]  = 1;
  ram[31061]  = 1;
  ram[31062]  = 1;
  ram[31063]  = 1;
  ram[31064]  = 1;
  ram[31065]  = 1;
  ram[31066]  = 1;
  ram[31067]  = 1;
  ram[31068]  = 1;
  ram[31069]  = 1;
  ram[31070]  = 1;
  ram[31071]  = 1;
  ram[31072]  = 1;
  ram[31073]  = 1;
  ram[31074]  = 1;
  ram[31075]  = 1;
  ram[31076]  = 1;
  ram[31077]  = 1;
  ram[31078]  = 1;
  ram[31079]  = 1;
  ram[31080]  = 1;
  ram[31081]  = 1;
  ram[31082]  = 1;
  ram[31083]  = 1;
  ram[31084]  = 1;
  ram[31085]  = 1;
  ram[31086]  = 1;
  ram[31087]  = 1;
  ram[31088]  = 1;
  ram[31089]  = 1;
  ram[31090]  = 1;
  ram[31091]  = 1;
  ram[31092]  = 1;
  ram[31093]  = 1;
  ram[31094]  = 1;
  ram[31095]  = 1;
  ram[31096]  = 1;
  ram[31097]  = 1;
  ram[31098]  = 1;
  ram[31099]  = 1;
  ram[31100]  = 1;
  ram[31101]  = 1;
  ram[31102]  = 1;
  ram[31103]  = 1;
  ram[31104]  = 1;
  ram[31105]  = 1;
  ram[31106]  = 1;
  ram[31107]  = 1;
  ram[31108]  = 1;
  ram[31109]  = 1;
  ram[31110]  = 1;
  ram[31111]  = 1;
  ram[31112]  = 1;
  ram[31113]  = 1;
  ram[31114]  = 1;
  ram[31115]  = 1;
  ram[31116]  = 1;
  ram[31117]  = 1;
  ram[31118]  = 1;
  ram[31119]  = 1;
  ram[31120]  = 1;
  ram[31121]  = 1;
  ram[31122]  = 1;
  ram[31123]  = 1;
  ram[31124]  = 1;
  ram[31125]  = 1;
  ram[31126]  = 1;
  ram[31127]  = 1;
  ram[31128]  = 1;
  ram[31129]  = 1;
  ram[31130]  = 1;
  ram[31131]  = 1;
  ram[31132]  = 1;
  ram[31133]  = 1;
  ram[31134]  = 1;
  ram[31135]  = 1;
  ram[31136]  = 1;
  ram[31137]  = 1;
  ram[31138]  = 1;
  ram[31139]  = 1;
  ram[31140]  = 1;
  ram[31141]  = 1;
  ram[31142]  = 1;
  ram[31143]  = 1;
  ram[31144]  = 1;
  ram[31145]  = 1;
  ram[31146]  = 1;
  ram[31147]  = 1;
  ram[31148]  = 1;
  ram[31149]  = 1;
  ram[31150]  = 1;
  ram[31151]  = 1;
  ram[31152]  = 1;
  ram[31153]  = 1;
  ram[31154]  = 1;
  ram[31155]  = 1;
  ram[31156]  = 1;
  ram[31157]  = 1;
  ram[31158]  = 1;
  ram[31159]  = 1;
  ram[31160]  = 1;
  ram[31161]  = 1;
  ram[31162]  = 1;
  ram[31163]  = 1;
  ram[31164]  = 1;
  ram[31165]  = 1;
  ram[31166]  = 1;
  ram[31167]  = 1;
  ram[31168]  = 1;
  ram[31169]  = 1;
  ram[31170]  = 1;
  ram[31171]  = 1;
  ram[31172]  = 1;
  ram[31173]  = 1;
  ram[31174]  = 1;
  ram[31175]  = 1;
  ram[31176]  = 1;
  ram[31177]  = 1;
  ram[31178]  = 1;
  ram[31179]  = 1;
  ram[31180]  = 1;
  ram[31181]  = 1;
  ram[31182]  = 1;
  ram[31183]  = 1;
  ram[31184]  = 1;
  ram[31185]  = 1;
  ram[31186]  = 1;
  ram[31187]  = 1;
  ram[31188]  = 1;
  ram[31189]  = 1;
  ram[31190]  = 1;
  ram[31191]  = 1;
  ram[31192]  = 1;
  ram[31193]  = 1;
  ram[31194]  = 1;
  ram[31195]  = 1;
  ram[31196]  = 1;
  ram[31197]  = 1;
  ram[31198]  = 1;
  ram[31199]  = 1;
  ram[31200]  = 1;
  ram[31201]  = 1;
  ram[31202]  = 1;
  ram[31203]  = 1;
  ram[31204]  = 1;
  ram[31205]  = 1;
  ram[31206]  = 1;
  ram[31207]  = 1;
  ram[31208]  = 1;
  ram[31209]  = 1;
  ram[31210]  = 1;
  ram[31211]  = 1;
  ram[31212]  = 1;
  ram[31213]  = 1;
  ram[31214]  = 1;
  ram[31215]  = 1;
  ram[31216]  = 1;
  ram[31217]  = 1;
  ram[31218]  = 1;
  ram[31219]  = 1;
  ram[31220]  = 1;
  ram[31221]  = 1;
  ram[31222]  = 1;
  ram[31223]  = 1;
  ram[31224]  = 1;
  ram[31225]  = 1;
  ram[31226]  = 1;
  ram[31227]  = 1;
  ram[31228]  = 1;
  ram[31229]  = 1;
  ram[31230]  = 1;
  ram[31231]  = 1;
  ram[31232]  = 1;
  ram[31233]  = 1;
  ram[31234]  = 1;
  ram[31235]  = 1;
  ram[31236]  = 1;
  ram[31237]  = 1;
  ram[31238]  = 1;
  ram[31239]  = 1;
  ram[31240]  = 1;
  ram[31241]  = 1;
  ram[31242]  = 1;
  ram[31243]  = 1;
  ram[31244]  = 1;
  ram[31245]  = 1;
  ram[31246]  = 1;
  ram[31247]  = 1;
  ram[31248]  = 1;
  ram[31249]  = 1;
  ram[31250]  = 1;
  ram[31251]  = 1;
  ram[31252]  = 1;
  ram[31253]  = 1;
  ram[31254]  = 1;
  ram[31255]  = 1;
  ram[31256]  = 1;
  ram[31257]  = 1;
  ram[31258]  = 0;
  ram[31259]  = 0;
  ram[31260]  = 1;
  ram[31261]  = 1;
  ram[31262]  = 1;
  ram[31263]  = 1;
  ram[31264]  = 1;
  ram[31265]  = 1;
  ram[31266]  = 1;
  ram[31267]  = 1;
  ram[31268]  = 1;
  ram[31269]  = 1;
  ram[31270]  = 1;
  ram[31271]  = 1;
  ram[31272]  = 1;
  ram[31273]  = 1;
  ram[31274]  = 1;
  ram[31275]  = 1;
  ram[31276]  = 1;
  ram[31277]  = 1;
  ram[31278]  = 1;
  ram[31279]  = 1;
  ram[31280]  = 1;
  ram[31281]  = 1;
  ram[31282]  = 1;
  ram[31283]  = 1;
  ram[31284]  = 1;
  ram[31285]  = 1;
  ram[31286]  = 1;
  ram[31287]  = 1;
  ram[31288]  = 1;
  ram[31289]  = 1;
  ram[31290]  = 1;
  ram[31291]  = 1;
  ram[31292]  = 1;
  ram[31293]  = 1;
  ram[31294]  = 1;
  ram[31295]  = 1;
  ram[31296]  = 1;
  ram[31297]  = 1;
  ram[31298]  = 1;
  ram[31299]  = 1;
  ram[31300]  = 1;
  ram[31301]  = 1;
  ram[31302]  = 1;
  ram[31303]  = 1;
  ram[31304]  = 1;
  ram[31305]  = 0;
  ram[31306]  = 0;
  ram[31307]  = 1;
  ram[31308]  = 1;
  ram[31309]  = 1;
  ram[31310]  = 1;
  ram[31311]  = 1;
  ram[31312]  = 1;
  ram[31313]  = 1;
  ram[31314]  = 1;
  ram[31315]  = 1;
  ram[31316]  = 1;
  ram[31317]  = 1;
  ram[31318]  = 1;
  ram[31319]  = 1;
  ram[31320]  = 1;
  ram[31321]  = 1;
  ram[31322]  = 1;
  ram[31323]  = 1;
  ram[31324]  = 1;
  ram[31325]  = 1;
  ram[31326]  = 1;
  ram[31327]  = 1;
  ram[31328]  = 1;
  ram[31329]  = 1;
  ram[31330]  = 0;
  ram[31331]  = 1;
  ram[31332]  = 1;
  ram[31333]  = 1;
  ram[31334]  = 1;
  ram[31335]  = 1;
  ram[31336]  = 1;
  ram[31337]  = 1;
  ram[31338]  = 1;
  ram[31339]  = 1;
  ram[31340]  = 1;
  ram[31341]  = 1;
  ram[31342]  = 1;
  ram[31343]  = 1;
  ram[31344]  = 1;
  ram[31345]  = 1;
  ram[31346]  = 1;
  ram[31347]  = 1;
  ram[31348]  = 1;
  ram[31349]  = 1;
  ram[31350]  = 1;
  ram[31351]  = 1;
  ram[31352]  = 1;
  ram[31353]  = 1;
  ram[31354]  = 1;
  ram[31355]  = 1;
  ram[31356]  = 1;
  ram[31357]  = 1;
  ram[31358]  = 1;
  ram[31359]  = 1;
  ram[31360]  = 1;
  ram[31361]  = 1;
  ram[31362]  = 1;
  ram[31363]  = 1;
  ram[31364]  = 1;
  ram[31365]  = 1;
  ram[31366]  = 1;
  ram[31367]  = 1;
  ram[31368]  = 1;
  ram[31369]  = 1;
  ram[31370]  = 1;
  ram[31371]  = 1;
  ram[31372]  = 1;
  ram[31373]  = 1;
  ram[31374]  = 1;
  ram[31375]  = 1;
  ram[31376]  = 1;
  ram[31377]  = 1;
  ram[31378]  = 1;
  ram[31379]  = 1;
  ram[31380]  = 1;
  ram[31381]  = 1;
  ram[31382]  = 1;
  ram[31383]  = 1;
  ram[31384]  = 1;
  ram[31385]  = 1;
  ram[31386]  = 1;
  ram[31387]  = 1;
  ram[31388]  = 1;
  ram[31389]  = 1;
  ram[31390]  = 1;
  ram[31391]  = 1;
  ram[31392]  = 1;
  ram[31393]  = 1;
  ram[31394]  = 1;
  ram[31395]  = 1;
  ram[31396]  = 1;
  ram[31397]  = 1;
  ram[31398]  = 1;
  ram[31399]  = 1;
  ram[31400]  = 1;
  ram[31401]  = 1;
  ram[31402]  = 1;
  ram[31403]  = 1;
  ram[31404]  = 1;
  ram[31405]  = 1;
  ram[31406]  = 1;
  ram[31407]  = 1;
  ram[31408]  = 1;
  ram[31409]  = 1;
  ram[31410]  = 1;
  ram[31411]  = 0;
  ram[31412]  = 1;
  ram[31413]  = 1;
  ram[31414]  = 1;
  ram[31415]  = 1;
  ram[31416]  = 1;
  ram[31417]  = 1;
  ram[31418]  = 1;
  ram[31419]  = 1;
  ram[31420]  = 1;
  ram[31421]  = 1;
  ram[31422]  = 1;
  ram[31423]  = 1;
  ram[31424]  = 1;
  ram[31425]  = 1;
  ram[31426]  = 1;
  ram[31427]  = 1;
  ram[31428]  = 1;
  ram[31429]  = 1;
  ram[31430]  = 1;
  ram[31431]  = 1;
  ram[31432]  = 1;
  ram[31433]  = 1;
  ram[31434]  = 1;
  ram[31435]  = 0;
  ram[31436]  = 0;
  ram[31437]  = 1;
  ram[31438]  = 1;
  ram[31439]  = 1;
  ram[31440]  = 1;
  ram[31441]  = 1;
  ram[31442]  = 1;
  ram[31443]  = 1;
  ram[31444]  = 1;
  ram[31445]  = 1;
  ram[31446]  = 1;
  ram[31447]  = 1;
  ram[31448]  = 1;
  ram[31449]  = 1;
  ram[31450]  = 1;
  ram[31451]  = 1;
  ram[31452]  = 1;
  ram[31453]  = 1;
  ram[31454]  = 1;
  ram[31455]  = 1;
  ram[31456]  = 1;
  ram[31457]  = 1;
  ram[31458]  = 1;
  ram[31459]  = 1;
  ram[31460]  = 1;
  ram[31461]  = 1;
  ram[31462]  = 1;
  ram[31463]  = 1;
  ram[31464]  = 1;
  ram[31465]  = 1;
  ram[31466]  = 1;
  ram[31467]  = 1;
  ram[31468]  = 1;
  ram[31469]  = 1;
  ram[31470]  = 1;
  ram[31471]  = 1;
  ram[31472]  = 1;
  ram[31473]  = 1;
  ram[31474]  = 1;
  ram[31475]  = 1;
  ram[31476]  = 1;
  ram[31477]  = 1;
  ram[31478]  = 1;
  ram[31479]  = 0;
  ram[31480]  = 1;
  ram[31481]  = 1;
  ram[31482]  = 1;
  ram[31483]  = 1;
  ram[31484]  = 1;
  ram[31485]  = 1;
  ram[31486]  = 1;
  ram[31487]  = 1;
  ram[31488]  = 1;
  ram[31489]  = 1;
  ram[31490]  = 1;
  ram[31491]  = 1;
  ram[31492]  = 1;
  ram[31493]  = 1;
  ram[31494]  = 1;
  ram[31495]  = 1;
  ram[31496]  = 1;
  ram[31497]  = 1;
  ram[31498]  = 1;
  ram[31499]  = 1;
  ram[31500]  = 1;
  ram[31501]  = 1;
  ram[31502]  = 1;
  ram[31503]  = 1;
  ram[31504]  = 1;
  ram[31505]  = 1;
  ram[31506]  = 1;
  ram[31507]  = 1;
  ram[31508]  = 1;
  ram[31509]  = 1;
  ram[31510]  = 1;
  ram[31511]  = 1;
  ram[31512]  = 1;
  ram[31513]  = 0;
  ram[31514]  = 1;
  ram[31515]  = 1;
  ram[31516]  = 1;
  ram[31517]  = 1;
  ram[31518]  = 1;
  ram[31519]  = 1;
  ram[31520]  = 1;
  ram[31521]  = 0;
  ram[31522]  = 1;
  ram[31523]  = 1;
  ram[31524]  = 1;
  ram[31525]  = 1;
  ram[31526]  = 1;
  ram[31527]  = 1;
  ram[31528]  = 1;
  ram[31529]  = 1;
  ram[31530]  = 1;
  ram[31531]  = 1;
  ram[31532]  = 1;
  ram[31533]  = 1;
  ram[31534]  = 1;
  ram[31535]  = 1;
  ram[31536]  = 1;
  ram[31537]  = 1;
  ram[31538]  = 1;
  ram[31539]  = 1;
  ram[31540]  = 1;
  ram[31541]  = 1;
  ram[31542]  = 1;
  ram[31543]  = 1;
  ram[31544]  = 1;
  ram[31545]  = 1;
  ram[31546]  = 1;
  ram[31547]  = 1;
  ram[31548]  = 1;
  ram[31549]  = 1;
  ram[31550]  = 1;
  ram[31551]  = 1;
  ram[31552]  = 1;
  ram[31553]  = 1;
  ram[31554]  = 1;
  ram[31555]  = 1;
  ram[31556]  = 1;
  ram[31557]  = 0;
  ram[31558]  = 0;
  ram[31559]  = 0;
  ram[31560]  = 0;
  ram[31561]  = 0;
  ram[31562]  = 1;
  ram[31563]  = 1;
  ram[31564]  = 1;
  ram[31565]  = 1;
  ram[31566]  = 1;
  ram[31567]  = 1;
  ram[31568]  = 1;
  ram[31569]  = 1;
  ram[31570]  = 1;
  ram[31571]  = 1;
  ram[31572]  = 1;
  ram[31573]  = 1;
  ram[31574]  = 1;
  ram[31575]  = 1;
  ram[31576]  = 1;
  ram[31577]  = 1;
  ram[31578]  = 1;
  ram[31579]  = 1;
  ram[31580]  = 1;
  ram[31581]  = 1;
  ram[31582]  = 1;
  ram[31583]  = 1;
  ram[31584]  = 1;
  ram[31585]  = 1;
  ram[31586]  = 1;
  ram[31587]  = 1;
  ram[31588]  = 1;
  ram[31589]  = 1;
  ram[31590]  = 1;
  ram[31591]  = 1;
  ram[31592]  = 1;
  ram[31593]  = 1;
  ram[31594]  = 1;
  ram[31595]  = 1;
  ram[31596]  = 1;
  ram[31597]  = 1;
  ram[31598]  = 1;
  ram[31599]  = 1;
  ram[31600]  = 1;
  ram[31601]  = 1;
  ram[31602]  = 1;
  ram[31603]  = 1;
  ram[31604]  = 1;
  ram[31605]  = 0;
  ram[31606]  = 0;
  ram[31607]  = 1;
  ram[31608]  = 1;
  ram[31609]  = 1;
  ram[31610]  = 1;
  ram[31611]  = 1;
  ram[31612]  = 1;
  ram[31613]  = 1;
  ram[31614]  = 1;
  ram[31615]  = 1;
  ram[31616]  = 1;
  ram[31617]  = 1;
  ram[31618]  = 1;
  ram[31619]  = 1;
  ram[31620]  = 1;
  ram[31621]  = 1;
  ram[31622]  = 1;
  ram[31623]  = 1;
  ram[31624]  = 1;
  ram[31625]  = 1;
  ram[31626]  = 1;
  ram[31627]  = 1;
  ram[31628]  = 1;
  ram[31629]  = 1;
  ram[31630]  = 0;
  ram[31631]  = 1;
  ram[31632]  = 1;
  ram[31633]  = 1;
  ram[31634]  = 1;
  ram[31635]  = 1;
  ram[31636]  = 1;
  ram[31637]  = 1;
  ram[31638]  = 1;
  ram[31639]  = 1;
  ram[31640]  = 1;
  ram[31641]  = 1;
  ram[31642]  = 1;
  ram[31643]  = 1;
  ram[31644]  = 1;
  ram[31645]  = 1;
  ram[31646]  = 1;
  ram[31647]  = 1;
  ram[31648]  = 1;
  ram[31649]  = 1;
  ram[31650]  = 1;
  ram[31651]  = 1;
  ram[31652]  = 1;
  ram[31653]  = 1;
  ram[31654]  = 1;
  ram[31655]  = 1;
  ram[31656]  = 1;
  ram[31657]  = 1;
  ram[31658]  = 1;
  ram[31659]  = 1;
  ram[31660]  = 1;
  ram[31661]  = 1;
  ram[31662]  = 1;
  ram[31663]  = 1;
  ram[31664]  = 1;
  ram[31665]  = 1;
  ram[31666]  = 1;
  ram[31667]  = 1;
  ram[31668]  = 1;
  ram[31669]  = 1;
  ram[31670]  = 1;
  ram[31671]  = 1;
  ram[31672]  = 1;
  ram[31673]  = 1;
  ram[31674]  = 1;
  ram[31675]  = 1;
  ram[31676]  = 1;
  ram[31677]  = 1;
  ram[31678]  = 1;
  ram[31679]  = 1;
  ram[31680]  = 1;
  ram[31681]  = 1;
  ram[31682]  = 1;
  ram[31683]  = 1;
  ram[31684]  = 1;
  ram[31685]  = 1;
  ram[31686]  = 1;
  ram[31687]  = 1;
  ram[31688]  = 1;
  ram[31689]  = 1;
  ram[31690]  = 1;
  ram[31691]  = 1;
  ram[31692]  = 1;
  ram[31693]  = 1;
  ram[31694]  = 1;
  ram[31695]  = 1;
  ram[31696]  = 1;
  ram[31697]  = 1;
  ram[31698]  = 1;
  ram[31699]  = 1;
  ram[31700]  = 1;
  ram[31701]  = 1;
  ram[31702]  = 1;
  ram[31703]  = 1;
  ram[31704]  = 1;
  ram[31705]  = 1;
  ram[31706]  = 1;
  ram[31707]  = 1;
  ram[31708]  = 1;
  ram[31709]  = 1;
  ram[31710]  = 1;
  ram[31711]  = 0;
  ram[31712]  = 1;
  ram[31713]  = 1;
  ram[31714]  = 1;
  ram[31715]  = 1;
  ram[31716]  = 1;
  ram[31717]  = 1;
  ram[31718]  = 1;
  ram[31719]  = 1;
  ram[31720]  = 1;
  ram[31721]  = 1;
  ram[31722]  = 1;
  ram[31723]  = 1;
  ram[31724]  = 1;
  ram[31725]  = 1;
  ram[31726]  = 1;
  ram[31727]  = 1;
  ram[31728]  = 1;
  ram[31729]  = 1;
  ram[31730]  = 1;
  ram[31731]  = 1;
  ram[31732]  = 1;
  ram[31733]  = 1;
  ram[31734]  = 1;
  ram[31735]  = 0;
  ram[31736]  = 0;
  ram[31737]  = 1;
  ram[31738]  = 1;
  ram[31739]  = 1;
  ram[31740]  = 1;
  ram[31741]  = 1;
  ram[31742]  = 1;
  ram[31743]  = 1;
  ram[31744]  = 1;
  ram[31745]  = 1;
  ram[31746]  = 1;
  ram[31747]  = 1;
  ram[31748]  = 1;
  ram[31749]  = 1;
  ram[31750]  = 1;
  ram[31751]  = 1;
  ram[31752]  = 1;
  ram[31753]  = 1;
  ram[31754]  = 1;
  ram[31755]  = 1;
  ram[31756]  = 1;
  ram[31757]  = 1;
  ram[31758]  = 1;
  ram[31759]  = 1;
  ram[31760]  = 1;
  ram[31761]  = 1;
  ram[31762]  = 1;
  ram[31763]  = 1;
  ram[31764]  = 1;
  ram[31765]  = 1;
  ram[31766]  = 1;
  ram[31767]  = 1;
  ram[31768]  = 1;
  ram[31769]  = 1;
  ram[31770]  = 1;
  ram[31771]  = 1;
  ram[31772]  = 1;
  ram[31773]  = 1;
  ram[31774]  = 1;
  ram[31775]  = 1;
  ram[31776]  = 1;
  ram[31777]  = 1;
  ram[31778]  = 1;
  ram[31779]  = 0;
  ram[31780]  = 1;
  ram[31781]  = 1;
  ram[31782]  = 1;
  ram[31783]  = 1;
  ram[31784]  = 1;
  ram[31785]  = 1;
  ram[31786]  = 1;
  ram[31787]  = 1;
  ram[31788]  = 1;
  ram[31789]  = 1;
  ram[31790]  = 1;
  ram[31791]  = 1;
  ram[31792]  = 1;
  ram[31793]  = 1;
  ram[31794]  = 1;
  ram[31795]  = 1;
  ram[31796]  = 1;
  ram[31797]  = 1;
  ram[31798]  = 1;
  ram[31799]  = 1;
  ram[31800]  = 1;
  ram[31801]  = 1;
  ram[31802]  = 1;
  ram[31803]  = 1;
  ram[31804]  = 1;
  ram[31805]  = 1;
  ram[31806]  = 1;
  ram[31807]  = 1;
  ram[31808]  = 1;
  ram[31809]  = 1;
  ram[31810]  = 1;
  ram[31811]  = 1;
  ram[31812]  = 1;
  ram[31813]  = 0;
  ram[31814]  = 1;
  ram[31815]  = 1;
  ram[31816]  = 1;
  ram[31817]  = 1;
  ram[31818]  = 1;
  ram[31819]  = 1;
  ram[31820]  = 0;
  ram[31821]  = 0;
  ram[31822]  = 1;
  ram[31823]  = 1;
  ram[31824]  = 1;
  ram[31825]  = 1;
  ram[31826]  = 1;
  ram[31827]  = 1;
  ram[31828]  = 1;
  ram[31829]  = 1;
  ram[31830]  = 1;
  ram[31831]  = 1;
  ram[31832]  = 1;
  ram[31833]  = 1;
  ram[31834]  = 1;
  ram[31835]  = 1;
  ram[31836]  = 1;
  ram[31837]  = 1;
  ram[31838]  = 1;
  ram[31839]  = 1;
  ram[31840]  = 1;
  ram[31841]  = 1;
  ram[31842]  = 1;
  ram[31843]  = 1;
  ram[31844]  = 1;
  ram[31845]  = 1;
  ram[31846]  = 1;
  ram[31847]  = 1;
  ram[31848]  = 1;
  ram[31849]  = 1;
  ram[31850]  = 1;
  ram[31851]  = 1;
  ram[31852]  = 1;
  ram[31853]  = 1;
  ram[31854]  = 1;
  ram[31855]  = 1;
  ram[31856]  = 0;
  ram[31857]  = 0;
  ram[31858]  = 1;
  ram[31859]  = 1;
  ram[31860]  = 0;
  ram[31861]  = 0;
  ram[31862]  = 1;
  ram[31863]  = 1;
  ram[31864]  = 1;
  ram[31865]  = 1;
  ram[31866]  = 1;
  ram[31867]  = 1;
  ram[31868]  = 1;
  ram[31869]  = 1;
  ram[31870]  = 1;
  ram[31871]  = 1;
  ram[31872]  = 1;
  ram[31873]  = 1;
  ram[31874]  = 1;
  ram[31875]  = 1;
  ram[31876]  = 1;
  ram[31877]  = 1;
  ram[31878]  = 1;
  ram[31879]  = 1;
  ram[31880]  = 1;
  ram[31881]  = 1;
  ram[31882]  = 1;
  ram[31883]  = 1;
  ram[31884]  = 1;
  ram[31885]  = 1;
  ram[31886]  = 1;
  ram[31887]  = 1;
  ram[31888]  = 1;
  ram[31889]  = 1;
  ram[31890]  = 1;
  ram[31891]  = 1;
  ram[31892]  = 1;
  ram[31893]  = 1;
  ram[31894]  = 1;
  ram[31895]  = 1;
  ram[31896]  = 1;
  ram[31897]  = 1;
  ram[31898]  = 1;
  ram[31899]  = 1;
  ram[31900]  = 1;
  ram[31901]  = 1;
  ram[31902]  = 1;
  ram[31903]  = 1;
  ram[31904]  = 1;
  ram[31905]  = 1;
  ram[31906]  = 1;
  ram[31907]  = 1;
  ram[31908]  = 1;
  ram[31909]  = 1;
  ram[31910]  = 1;
  ram[31911]  = 1;
  ram[31912]  = 1;
  ram[31913]  = 1;
  ram[31914]  = 1;
  ram[31915]  = 1;
  ram[31916]  = 1;
  ram[31917]  = 1;
  ram[31918]  = 1;
  ram[31919]  = 1;
  ram[31920]  = 1;
  ram[31921]  = 1;
  ram[31922]  = 1;
  ram[31923]  = 1;
  ram[31924]  = 1;
  ram[31925]  = 1;
  ram[31926]  = 1;
  ram[31927]  = 1;
  ram[31928]  = 1;
  ram[31929]  = 1;
  ram[31930]  = 0;
  ram[31931]  = 1;
  ram[31932]  = 1;
  ram[31933]  = 1;
  ram[31934]  = 1;
  ram[31935]  = 1;
  ram[31936]  = 1;
  ram[31937]  = 1;
  ram[31938]  = 1;
  ram[31939]  = 1;
  ram[31940]  = 1;
  ram[31941]  = 1;
  ram[31942]  = 1;
  ram[31943]  = 1;
  ram[31944]  = 1;
  ram[31945]  = 1;
  ram[31946]  = 1;
  ram[31947]  = 1;
  ram[31948]  = 1;
  ram[31949]  = 1;
  ram[31950]  = 1;
  ram[31951]  = 1;
  ram[31952]  = 1;
  ram[31953]  = 1;
  ram[31954]  = 1;
  ram[31955]  = 1;
  ram[31956]  = 1;
  ram[31957]  = 1;
  ram[31958]  = 1;
  ram[31959]  = 1;
  ram[31960]  = 1;
  ram[31961]  = 1;
  ram[31962]  = 1;
  ram[31963]  = 1;
  ram[31964]  = 1;
  ram[31965]  = 1;
  ram[31966]  = 1;
  ram[31967]  = 1;
  ram[31968]  = 1;
  ram[31969]  = 1;
  ram[31970]  = 1;
  ram[31971]  = 1;
  ram[31972]  = 1;
  ram[31973]  = 1;
  ram[31974]  = 1;
  ram[31975]  = 1;
  ram[31976]  = 1;
  ram[31977]  = 1;
  ram[31978]  = 1;
  ram[31979]  = 1;
  ram[31980]  = 1;
  ram[31981]  = 1;
  ram[31982]  = 1;
  ram[31983]  = 1;
  ram[31984]  = 1;
  ram[31985]  = 1;
  ram[31986]  = 1;
  ram[31987]  = 1;
  ram[31988]  = 1;
  ram[31989]  = 1;
  ram[31990]  = 1;
  ram[31991]  = 1;
  ram[31992]  = 1;
  ram[31993]  = 1;
  ram[31994]  = 1;
  ram[31995]  = 1;
  ram[31996]  = 1;
  ram[31997]  = 1;
  ram[31998]  = 1;
  ram[31999]  = 1;
  ram[32000]  = 1;
  ram[32001]  = 1;
  ram[32002]  = 1;
  ram[32003]  = 1;
  ram[32004]  = 1;
  ram[32005]  = 1;
  ram[32006]  = 1;
  ram[32007]  = 1;
  ram[32008]  = 1;
  ram[32009]  = 1;
  ram[32010]  = 1;
  ram[32011]  = 0;
  ram[32012]  = 1;
  ram[32013]  = 1;
  ram[32014]  = 1;
  ram[32015]  = 1;
  ram[32016]  = 1;
  ram[32017]  = 1;
  ram[32018]  = 1;
  ram[32019]  = 1;
  ram[32020]  = 1;
  ram[32021]  = 1;
  ram[32022]  = 1;
  ram[32023]  = 1;
  ram[32024]  = 1;
  ram[32025]  = 1;
  ram[32026]  = 1;
  ram[32027]  = 1;
  ram[32028]  = 1;
  ram[32029]  = 1;
  ram[32030]  = 1;
  ram[32031]  = 1;
  ram[32032]  = 1;
  ram[32033]  = 1;
  ram[32034]  = 1;
  ram[32035]  = 0;
  ram[32036]  = 0;
  ram[32037]  = 1;
  ram[32038]  = 1;
  ram[32039]  = 1;
  ram[32040]  = 1;
  ram[32041]  = 1;
  ram[32042]  = 1;
  ram[32043]  = 1;
  ram[32044]  = 1;
  ram[32045]  = 1;
  ram[32046]  = 1;
  ram[32047]  = 1;
  ram[32048]  = 1;
  ram[32049]  = 1;
  ram[32050]  = 1;
  ram[32051]  = 1;
  ram[32052]  = 1;
  ram[32053]  = 1;
  ram[32054]  = 1;
  ram[32055]  = 1;
  ram[32056]  = 1;
  ram[32057]  = 1;
  ram[32058]  = 1;
  ram[32059]  = 1;
  ram[32060]  = 1;
  ram[32061]  = 1;
  ram[32062]  = 1;
  ram[32063]  = 1;
  ram[32064]  = 1;
  ram[32065]  = 1;
  ram[32066]  = 1;
  ram[32067]  = 1;
  ram[32068]  = 1;
  ram[32069]  = 1;
  ram[32070]  = 1;
  ram[32071]  = 1;
  ram[32072]  = 1;
  ram[32073]  = 1;
  ram[32074]  = 1;
  ram[32075]  = 1;
  ram[32076]  = 1;
  ram[32077]  = 1;
  ram[32078]  = 1;
  ram[32079]  = 0;
  ram[32080]  = 1;
  ram[32081]  = 1;
  ram[32082]  = 1;
  ram[32083]  = 1;
  ram[32084]  = 1;
  ram[32085]  = 1;
  ram[32086]  = 1;
  ram[32087]  = 1;
  ram[32088]  = 1;
  ram[32089]  = 1;
  ram[32090]  = 1;
  ram[32091]  = 1;
  ram[32092]  = 1;
  ram[32093]  = 1;
  ram[32094]  = 1;
  ram[32095]  = 1;
  ram[32096]  = 1;
  ram[32097]  = 1;
  ram[32098]  = 1;
  ram[32099]  = 1;
  ram[32100]  = 1;
  ram[32101]  = 1;
  ram[32102]  = 1;
  ram[32103]  = 1;
  ram[32104]  = 1;
  ram[32105]  = 1;
  ram[32106]  = 1;
  ram[32107]  = 1;
  ram[32108]  = 1;
  ram[32109]  = 1;
  ram[32110]  = 1;
  ram[32111]  = 1;
  ram[32112]  = 1;
  ram[32113]  = 0;
  ram[32114]  = 0;
  ram[32115]  = 1;
  ram[32116]  = 1;
  ram[32117]  = 1;
  ram[32118]  = 1;
  ram[32119]  = 1;
  ram[32120]  = 0;
  ram[32121]  = 1;
  ram[32122]  = 1;
  ram[32123]  = 1;
  ram[32124]  = 1;
  ram[32125]  = 1;
  ram[32126]  = 1;
  ram[32127]  = 1;
  ram[32128]  = 1;
  ram[32129]  = 1;
  ram[32130]  = 1;
  ram[32131]  = 1;
  ram[32132]  = 1;
  ram[32133]  = 1;
  ram[32134]  = 1;
  ram[32135]  = 1;
  ram[32136]  = 1;
  ram[32137]  = 1;
  ram[32138]  = 1;
  ram[32139]  = 1;
  ram[32140]  = 1;
  ram[32141]  = 1;
  ram[32142]  = 1;
  ram[32143]  = 1;
  ram[32144]  = 1;
  ram[32145]  = 1;
  ram[32146]  = 1;
  ram[32147]  = 1;
  ram[32148]  = 1;
  ram[32149]  = 1;
  ram[32150]  = 1;
  ram[32151]  = 1;
  ram[32152]  = 1;
  ram[32153]  = 1;
  ram[32154]  = 1;
  ram[32155]  = 1;
  ram[32156]  = 0;
  ram[32157]  = 1;
  ram[32158]  = 1;
  ram[32159]  = 1;
  ram[32160]  = 1;
  ram[32161]  = 0;
  ram[32162]  = 0;
  ram[32163]  = 1;
  ram[32164]  = 1;
  ram[32165]  = 1;
  ram[32166]  = 1;
  ram[32167]  = 1;
  ram[32168]  = 1;
  ram[32169]  = 1;
  ram[32170]  = 1;
  ram[32171]  = 1;
  ram[32172]  = 1;
  ram[32173]  = 1;
  ram[32174]  = 1;
  ram[32175]  = 1;
  ram[32176]  = 1;
  ram[32177]  = 1;
  ram[32178]  = 1;
  ram[32179]  = 1;
  ram[32180]  = 1;
  ram[32181]  = 1;
  ram[32182]  = 1;
  ram[32183]  = 1;
  ram[32184]  = 1;
  ram[32185]  = 1;
  ram[32186]  = 1;
  ram[32187]  = 1;
  ram[32188]  = 1;
  ram[32189]  = 1;
  ram[32190]  = 1;
  ram[32191]  = 1;
  ram[32192]  = 1;
  ram[32193]  = 1;
  ram[32194]  = 1;
  ram[32195]  = 1;
  ram[32196]  = 1;
  ram[32197]  = 1;
  ram[32198]  = 1;
  ram[32199]  = 1;
  ram[32200]  = 1;
  ram[32201]  = 1;
  ram[32202]  = 1;
  ram[32203]  = 1;
  ram[32204]  = 1;
  ram[32205]  = 1;
  ram[32206]  = 1;
  ram[32207]  = 1;
  ram[32208]  = 1;
  ram[32209]  = 1;
  ram[32210]  = 1;
  ram[32211]  = 1;
  ram[32212]  = 1;
  ram[32213]  = 1;
  ram[32214]  = 1;
  ram[32215]  = 1;
  ram[32216]  = 1;
  ram[32217]  = 1;
  ram[32218]  = 1;
  ram[32219]  = 1;
  ram[32220]  = 1;
  ram[32221]  = 1;
  ram[32222]  = 1;
  ram[32223]  = 1;
  ram[32224]  = 1;
  ram[32225]  = 1;
  ram[32226]  = 1;
  ram[32227]  = 1;
  ram[32228]  = 1;
  ram[32229]  = 1;
  ram[32230]  = 0;
  ram[32231]  = 1;
  ram[32232]  = 1;
  ram[32233]  = 1;
  ram[32234]  = 1;
  ram[32235]  = 1;
  ram[32236]  = 1;
  ram[32237]  = 1;
  ram[32238]  = 1;
  ram[32239]  = 1;
  ram[32240]  = 1;
  ram[32241]  = 1;
  ram[32242]  = 1;
  ram[32243]  = 1;
  ram[32244]  = 1;
  ram[32245]  = 1;
  ram[32246]  = 1;
  ram[32247]  = 1;
  ram[32248]  = 1;
  ram[32249]  = 1;
  ram[32250]  = 1;
  ram[32251]  = 1;
  ram[32252]  = 1;
  ram[32253]  = 1;
  ram[32254]  = 1;
  ram[32255]  = 1;
  ram[32256]  = 1;
  ram[32257]  = 1;
  ram[32258]  = 1;
  ram[32259]  = 1;
  ram[32260]  = 1;
  ram[32261]  = 1;
  ram[32262]  = 1;
  ram[32263]  = 1;
  ram[32264]  = 1;
  ram[32265]  = 1;
  ram[32266]  = 1;
  ram[32267]  = 1;
  ram[32268]  = 1;
  ram[32269]  = 1;
  ram[32270]  = 1;
  ram[32271]  = 1;
  ram[32272]  = 1;
  ram[32273]  = 1;
  ram[32274]  = 1;
  ram[32275]  = 1;
  ram[32276]  = 1;
  ram[32277]  = 1;
  ram[32278]  = 1;
  ram[32279]  = 1;
  ram[32280]  = 1;
  ram[32281]  = 1;
  ram[32282]  = 1;
  ram[32283]  = 1;
  ram[32284]  = 1;
  ram[32285]  = 1;
  ram[32286]  = 1;
  ram[32287]  = 1;
  ram[32288]  = 1;
  ram[32289]  = 1;
  ram[32290]  = 1;
  ram[32291]  = 1;
  ram[32292]  = 1;
  ram[32293]  = 1;
  ram[32294]  = 1;
  ram[32295]  = 1;
  ram[32296]  = 1;
  ram[32297]  = 1;
  ram[32298]  = 1;
  ram[32299]  = 1;
  ram[32300]  = 1;
  ram[32301]  = 1;
  ram[32302]  = 1;
  ram[32303]  = 1;
  ram[32304]  = 1;
  ram[32305]  = 0;
  ram[32306]  = 1;
  ram[32307]  = 1;
  ram[32308]  = 1;
  ram[32309]  = 1;
  ram[32310]  = 1;
  ram[32311]  = 0;
  ram[32312]  = 1;
  ram[32313]  = 1;
  ram[32314]  = 1;
  ram[32315]  = 1;
  ram[32316]  = 1;
  ram[32317]  = 1;
  ram[32318]  = 1;
  ram[32319]  = 1;
  ram[32320]  = 1;
  ram[32321]  = 1;
  ram[32322]  = 1;
  ram[32323]  = 1;
  ram[32324]  = 1;
  ram[32325]  = 1;
  ram[32326]  = 1;
  ram[32327]  = 1;
  ram[32328]  = 1;
  ram[32329]  = 1;
  ram[32330]  = 1;
  ram[32331]  = 1;
  ram[32332]  = 1;
  ram[32333]  = 1;
  ram[32334]  = 1;
  ram[32335]  = 0;
  ram[32336]  = 0;
  ram[32337]  = 1;
  ram[32338]  = 1;
  ram[32339]  = 1;
  ram[32340]  = 1;
  ram[32341]  = 1;
  ram[32342]  = 1;
  ram[32343]  = 1;
  ram[32344]  = 1;
  ram[32345]  = 1;
  ram[32346]  = 1;
  ram[32347]  = 1;
  ram[32348]  = 1;
  ram[32349]  = 1;
  ram[32350]  = 1;
  ram[32351]  = 1;
  ram[32352]  = 1;
  ram[32353]  = 1;
  ram[32354]  = 1;
  ram[32355]  = 1;
  ram[32356]  = 1;
  ram[32357]  = 1;
  ram[32358]  = 1;
  ram[32359]  = 1;
  ram[32360]  = 1;
  ram[32361]  = 1;
  ram[32362]  = 1;
  ram[32363]  = 1;
  ram[32364]  = 1;
  ram[32365]  = 1;
  ram[32366]  = 1;
  ram[32367]  = 1;
  ram[32368]  = 1;
  ram[32369]  = 1;
  ram[32370]  = 1;
  ram[32371]  = 1;
  ram[32372]  = 1;
  ram[32373]  = 1;
  ram[32374]  = 1;
  ram[32375]  = 1;
  ram[32376]  = 1;
  ram[32377]  = 1;
  ram[32378]  = 1;
  ram[32379]  = 0;
  ram[32380]  = 1;
  ram[32381]  = 1;
  ram[32382]  = 1;
  ram[32383]  = 1;
  ram[32384]  = 1;
  ram[32385]  = 1;
  ram[32386]  = 1;
  ram[32387]  = 1;
  ram[32388]  = 1;
  ram[32389]  = 1;
  ram[32390]  = 1;
  ram[32391]  = 1;
  ram[32392]  = 1;
  ram[32393]  = 1;
  ram[32394]  = 1;
  ram[32395]  = 1;
  ram[32396]  = 1;
  ram[32397]  = 1;
  ram[32398]  = 1;
  ram[32399]  = 1;
  ram[32400]  = 1;
  ram[32401]  = 1;
  ram[32402]  = 1;
  ram[32403]  = 1;
  ram[32404]  = 1;
  ram[32405]  = 1;
  ram[32406]  = 1;
  ram[32407]  = 1;
  ram[32408]  = 1;
  ram[32409]  = 1;
  ram[32410]  = 1;
  ram[32411]  = 1;
  ram[32412]  = 1;
  ram[32413]  = 1;
  ram[32414]  = 0;
  ram[32415]  = 1;
  ram[32416]  = 1;
  ram[32417]  = 1;
  ram[32418]  = 1;
  ram[32419]  = 1;
  ram[32420]  = 0;
  ram[32421]  = 1;
  ram[32422]  = 1;
  ram[32423]  = 1;
  ram[32424]  = 1;
  ram[32425]  = 1;
  ram[32426]  = 1;
  ram[32427]  = 1;
  ram[32428]  = 1;
  ram[32429]  = 1;
  ram[32430]  = 1;
  ram[32431]  = 1;
  ram[32432]  = 1;
  ram[32433]  = 1;
  ram[32434]  = 1;
  ram[32435]  = 1;
  ram[32436]  = 1;
  ram[32437]  = 1;
  ram[32438]  = 1;
  ram[32439]  = 1;
  ram[32440]  = 1;
  ram[32441]  = 1;
  ram[32442]  = 1;
  ram[32443]  = 1;
  ram[32444]  = 1;
  ram[32445]  = 1;
  ram[32446]  = 1;
  ram[32447]  = 1;
  ram[32448]  = 1;
  ram[32449]  = 1;
  ram[32450]  = 1;
  ram[32451]  = 1;
  ram[32452]  = 1;
  ram[32453]  = 1;
  ram[32454]  = 1;
  ram[32455]  = 1;
  ram[32456]  = 0;
  ram[32457]  = 1;
  ram[32458]  = 1;
  ram[32459]  = 1;
  ram[32460]  = 1;
  ram[32461]  = 1;
  ram[32462]  = 0;
  ram[32463]  = 1;
  ram[32464]  = 1;
  ram[32465]  = 1;
  ram[32466]  = 1;
  ram[32467]  = 1;
  ram[32468]  = 1;
  ram[32469]  = 1;
  ram[32470]  = 1;
  ram[32471]  = 1;
  ram[32472]  = 1;
  ram[32473]  = 1;
  ram[32474]  = 1;
  ram[32475]  = 1;
  ram[32476]  = 1;
  ram[32477]  = 1;
  ram[32478]  = 1;
  ram[32479]  = 1;
  ram[32480]  = 1;
  ram[32481]  = 1;
  ram[32482]  = 1;
  ram[32483]  = 1;
  ram[32484]  = 1;
  ram[32485]  = 1;
  ram[32486]  = 1;
  ram[32487]  = 1;
  ram[32488]  = 1;
  ram[32489]  = 1;
  ram[32490]  = 1;
  ram[32491]  = 1;
  ram[32492]  = 1;
  ram[32493]  = 1;
  ram[32494]  = 1;
  ram[32495]  = 1;
  ram[32496]  = 1;
  ram[32497]  = 1;
  ram[32498]  = 1;
  ram[32499]  = 1;
  ram[32500]  = 1;
  ram[32501]  = 1;
  ram[32502]  = 1;
  ram[32503]  = 1;
  ram[32504]  = 1;
  ram[32505]  = 1;
  ram[32506]  = 1;
  ram[32507]  = 1;
  ram[32508]  = 1;
  ram[32509]  = 1;
  ram[32510]  = 1;
  ram[32511]  = 1;
  ram[32512]  = 1;
  ram[32513]  = 1;
  ram[32514]  = 1;
  ram[32515]  = 1;
  ram[32516]  = 1;
  ram[32517]  = 1;
  ram[32518]  = 1;
  ram[32519]  = 1;
  ram[32520]  = 1;
  ram[32521]  = 1;
  ram[32522]  = 1;
  ram[32523]  = 1;
  ram[32524]  = 1;
  ram[32525]  = 1;
  ram[32526]  = 1;
  ram[32527]  = 1;
  ram[32528]  = 1;
  ram[32529]  = 1;
  ram[32530]  = 0;
  ram[32531]  = 1;
  ram[32532]  = 1;
  ram[32533]  = 1;
  ram[32534]  = 1;
  ram[32535]  = 1;
  ram[32536]  = 1;
  ram[32537]  = 1;
  ram[32538]  = 1;
  ram[32539]  = 1;
  ram[32540]  = 1;
  ram[32541]  = 1;
  ram[32542]  = 1;
  ram[32543]  = 1;
  ram[32544]  = 1;
  ram[32545]  = 1;
  ram[32546]  = 1;
  ram[32547]  = 1;
  ram[32548]  = 1;
  ram[32549]  = 1;
  ram[32550]  = 1;
  ram[32551]  = 1;
  ram[32552]  = 1;
  ram[32553]  = 1;
  ram[32554]  = 1;
  ram[32555]  = 1;
  ram[32556]  = 1;
  ram[32557]  = 1;
  ram[32558]  = 1;
  ram[32559]  = 1;
  ram[32560]  = 1;
  ram[32561]  = 1;
  ram[32562]  = 1;
  ram[32563]  = 1;
  ram[32564]  = 1;
  ram[32565]  = 1;
  ram[32566]  = 1;
  ram[32567]  = 1;
  ram[32568]  = 1;
  ram[32569]  = 1;
  ram[32570]  = 1;
  ram[32571]  = 1;
  ram[32572]  = 1;
  ram[32573]  = 1;
  ram[32574]  = 1;
  ram[32575]  = 1;
  ram[32576]  = 1;
  ram[32577]  = 1;
  ram[32578]  = 1;
  ram[32579]  = 1;
  ram[32580]  = 1;
  ram[32581]  = 1;
  ram[32582]  = 1;
  ram[32583]  = 1;
  ram[32584]  = 1;
  ram[32585]  = 1;
  ram[32586]  = 1;
  ram[32587]  = 1;
  ram[32588]  = 1;
  ram[32589]  = 1;
  ram[32590]  = 1;
  ram[32591]  = 1;
  ram[32592]  = 1;
  ram[32593]  = 1;
  ram[32594]  = 1;
  ram[32595]  = 1;
  ram[32596]  = 1;
  ram[32597]  = 1;
  ram[32598]  = 1;
  ram[32599]  = 1;
  ram[32600]  = 1;
  ram[32601]  = 1;
  ram[32602]  = 1;
  ram[32603]  = 1;
  ram[32604]  = 1;
  ram[32605]  = 0;
  ram[32606]  = 1;
  ram[32607]  = 1;
  ram[32608]  = 1;
  ram[32609]  = 1;
  ram[32610]  = 1;
  ram[32611]  = 0;
  ram[32612]  = 1;
  ram[32613]  = 1;
  ram[32614]  = 1;
  ram[32615]  = 1;
  ram[32616]  = 1;
  ram[32617]  = 1;
  ram[32618]  = 1;
  ram[32619]  = 1;
  ram[32620]  = 1;
  ram[32621]  = 1;
  ram[32622]  = 1;
  ram[32623]  = 1;
  ram[32624]  = 1;
  ram[32625]  = 1;
  ram[32626]  = 1;
  ram[32627]  = 1;
  ram[32628]  = 1;
  ram[32629]  = 1;
  ram[32630]  = 1;
  ram[32631]  = 1;
  ram[32632]  = 1;
  ram[32633]  = 1;
  ram[32634]  = 1;
  ram[32635]  = 0;
  ram[32636]  = 0;
  ram[32637]  = 1;
  ram[32638]  = 1;
  ram[32639]  = 1;
  ram[32640]  = 1;
  ram[32641]  = 1;
  ram[32642]  = 1;
  ram[32643]  = 1;
  ram[32644]  = 1;
  ram[32645]  = 1;
  ram[32646]  = 1;
  ram[32647]  = 1;
  ram[32648]  = 1;
  ram[32649]  = 1;
  ram[32650]  = 1;
  ram[32651]  = 1;
  ram[32652]  = 1;
  ram[32653]  = 1;
  ram[32654]  = 1;
  ram[32655]  = 1;
  ram[32656]  = 1;
  ram[32657]  = 1;
  ram[32658]  = 1;
  ram[32659]  = 1;
  ram[32660]  = 1;
  ram[32661]  = 1;
  ram[32662]  = 1;
  ram[32663]  = 1;
  ram[32664]  = 1;
  ram[32665]  = 1;
  ram[32666]  = 1;
  ram[32667]  = 1;
  ram[32668]  = 1;
  ram[32669]  = 1;
  ram[32670]  = 1;
  ram[32671]  = 1;
  ram[32672]  = 1;
  ram[32673]  = 1;
  ram[32674]  = 1;
  ram[32675]  = 1;
  ram[32676]  = 1;
  ram[32677]  = 1;
  ram[32678]  = 1;
  ram[32679]  = 0;
  ram[32680]  = 1;
  ram[32681]  = 1;
  ram[32682]  = 1;
  ram[32683]  = 1;
  ram[32684]  = 1;
  ram[32685]  = 1;
  ram[32686]  = 1;
  ram[32687]  = 1;
  ram[32688]  = 1;
  ram[32689]  = 1;
  ram[32690]  = 1;
  ram[32691]  = 1;
  ram[32692]  = 1;
  ram[32693]  = 1;
  ram[32694]  = 1;
  ram[32695]  = 1;
  ram[32696]  = 1;
  ram[32697]  = 1;
  ram[32698]  = 1;
  ram[32699]  = 1;
  ram[32700]  = 1;
  ram[32701]  = 1;
  ram[32702]  = 1;
  ram[32703]  = 1;
  ram[32704]  = 1;
  ram[32705]  = 1;
  ram[32706]  = 1;
  ram[32707]  = 1;
  ram[32708]  = 1;
  ram[32709]  = 1;
  ram[32710]  = 1;
  ram[32711]  = 1;
  ram[32712]  = 1;
  ram[32713]  = 1;
  ram[32714]  = 0;
  ram[32715]  = 1;
  ram[32716]  = 1;
  ram[32717]  = 1;
  ram[32718]  = 1;
  ram[32719]  = 0;
  ram[32720]  = 0;
  ram[32721]  = 1;
  ram[32722]  = 1;
  ram[32723]  = 1;
  ram[32724]  = 1;
  ram[32725]  = 1;
  ram[32726]  = 1;
  ram[32727]  = 1;
  ram[32728]  = 1;
  ram[32729]  = 1;
  ram[32730]  = 1;
  ram[32731]  = 1;
  ram[32732]  = 1;
  ram[32733]  = 1;
  ram[32734]  = 1;
  ram[32735]  = 1;
  ram[32736]  = 1;
  ram[32737]  = 1;
  ram[32738]  = 1;
  ram[32739]  = 1;
  ram[32740]  = 1;
  ram[32741]  = 1;
  ram[32742]  = 1;
  ram[32743]  = 1;
  ram[32744]  = 1;
  ram[32745]  = 1;
  ram[32746]  = 1;
  ram[32747]  = 1;
  ram[32748]  = 1;
  ram[32749]  = 1;
  ram[32750]  = 1;
  ram[32751]  = 1;
  ram[32752]  = 1;
  ram[32753]  = 1;
  ram[32754]  = 1;
  ram[32755]  = 1;
  ram[32756]  = 0;
  ram[32757]  = 1;
  ram[32758]  = 1;
  ram[32759]  = 1;
  ram[32760]  = 1;
  ram[32761]  = 1;
  ram[32762]  = 0;
  ram[32763]  = 1;
  ram[32764]  = 1;
  ram[32765]  = 1;
  ram[32766]  = 1;
  ram[32767]  = 1;
  ram[32768]  = 1;
  ram[32769]  = 1;
  ram[32770]  = 1;
  ram[32771]  = 1;
  ram[32772]  = 1;
  ram[32773]  = 1;
  ram[32774]  = 1;
  ram[32775]  = 1;
  ram[32776]  = 1;
  ram[32777]  = 1;
  ram[32778]  = 1;
  ram[32779]  = 1;
  ram[32780]  = 1;
  ram[32781]  = 1;
  ram[32782]  = 1;
  ram[32783]  = 1;
  ram[32784]  = 1;
  ram[32785]  = 1;
  ram[32786]  = 1;
  ram[32787]  = 1;
  ram[32788]  = 1;
  ram[32789]  = 1;
  ram[32790]  = 1;
  ram[32791]  = 1;
  ram[32792]  = 1;
  ram[32793]  = 1;
  ram[32794]  = 1;
  ram[32795]  = 1;
  ram[32796]  = 1;
  ram[32797]  = 1;
  ram[32798]  = 1;
  ram[32799]  = 1;
  ram[32800]  = 1;
  ram[32801]  = 1;
  ram[32802]  = 1;
  ram[32803]  = 1;
  ram[32804]  = 1;
  ram[32805]  = 1;
  ram[32806]  = 1;
  ram[32807]  = 1;
  ram[32808]  = 1;
  ram[32809]  = 1;
  ram[32810]  = 1;
  ram[32811]  = 1;
  ram[32812]  = 1;
  ram[32813]  = 1;
  ram[32814]  = 1;
  ram[32815]  = 1;
  ram[32816]  = 1;
  ram[32817]  = 1;
  ram[32818]  = 1;
  ram[32819]  = 1;
  ram[32820]  = 1;
  ram[32821]  = 1;
  ram[32822]  = 1;
  ram[32823]  = 1;
  ram[32824]  = 1;
  ram[32825]  = 1;
  ram[32826]  = 1;
  ram[32827]  = 1;
  ram[32828]  = 1;
  ram[32829]  = 1;
  ram[32830]  = 0;
  ram[32831]  = 1;
  ram[32832]  = 1;
  ram[32833]  = 1;
  ram[32834]  = 1;
  ram[32835]  = 1;
  ram[32836]  = 1;
  ram[32837]  = 1;
  ram[32838]  = 1;
  ram[32839]  = 1;
  ram[32840]  = 1;
  ram[32841]  = 1;
  ram[32842]  = 1;
  ram[32843]  = 1;
  ram[32844]  = 1;
  ram[32845]  = 1;
  ram[32846]  = 1;
  ram[32847]  = 1;
  ram[32848]  = 1;
  ram[32849]  = 1;
  ram[32850]  = 1;
  ram[32851]  = 1;
  ram[32852]  = 1;
  ram[32853]  = 1;
  ram[32854]  = 1;
  ram[32855]  = 1;
  ram[32856]  = 1;
  ram[32857]  = 1;
  ram[32858]  = 1;
  ram[32859]  = 1;
  ram[32860]  = 1;
  ram[32861]  = 1;
  ram[32862]  = 1;
  ram[32863]  = 1;
  ram[32864]  = 1;
  ram[32865]  = 1;
  ram[32866]  = 1;
  ram[32867]  = 1;
  ram[32868]  = 1;
  ram[32869]  = 1;
  ram[32870]  = 1;
  ram[32871]  = 1;
  ram[32872]  = 1;
  ram[32873]  = 1;
  ram[32874]  = 1;
  ram[32875]  = 1;
  ram[32876]  = 1;
  ram[32877]  = 1;
  ram[32878]  = 1;
  ram[32879]  = 1;
  ram[32880]  = 1;
  ram[32881]  = 1;
  ram[32882]  = 1;
  ram[32883]  = 1;
  ram[32884]  = 1;
  ram[32885]  = 1;
  ram[32886]  = 1;
  ram[32887]  = 1;
  ram[32888]  = 1;
  ram[32889]  = 1;
  ram[32890]  = 1;
  ram[32891]  = 1;
  ram[32892]  = 1;
  ram[32893]  = 1;
  ram[32894]  = 1;
  ram[32895]  = 1;
  ram[32896]  = 1;
  ram[32897]  = 1;
  ram[32898]  = 1;
  ram[32899]  = 1;
  ram[32900]  = 1;
  ram[32901]  = 1;
  ram[32902]  = 1;
  ram[32903]  = 1;
  ram[32904]  = 1;
  ram[32905]  = 0;
  ram[32906]  = 1;
  ram[32907]  = 1;
  ram[32908]  = 1;
  ram[32909]  = 1;
  ram[32910]  = 1;
  ram[32911]  = 0;
  ram[32912]  = 1;
  ram[32913]  = 1;
  ram[32914]  = 1;
  ram[32915]  = 1;
  ram[32916]  = 1;
  ram[32917]  = 1;
  ram[32918]  = 1;
  ram[32919]  = 1;
  ram[32920]  = 1;
  ram[32921]  = 1;
  ram[32922]  = 1;
  ram[32923]  = 1;
  ram[32924]  = 1;
  ram[32925]  = 1;
  ram[32926]  = 1;
  ram[32927]  = 1;
  ram[32928]  = 1;
  ram[32929]  = 1;
  ram[32930]  = 1;
  ram[32931]  = 1;
  ram[32932]  = 1;
  ram[32933]  = 1;
  ram[32934]  = 1;
  ram[32935]  = 0;
  ram[32936]  = 0;
  ram[32937]  = 1;
  ram[32938]  = 1;
  ram[32939]  = 1;
  ram[32940]  = 1;
  ram[32941]  = 1;
  ram[32942]  = 1;
  ram[32943]  = 1;
  ram[32944]  = 1;
  ram[32945]  = 1;
  ram[32946]  = 1;
  ram[32947]  = 1;
  ram[32948]  = 1;
  ram[32949]  = 1;
  ram[32950]  = 1;
  ram[32951]  = 1;
  ram[32952]  = 1;
  ram[32953]  = 1;
  ram[32954]  = 1;
  ram[32955]  = 1;
  ram[32956]  = 1;
  ram[32957]  = 1;
  ram[32958]  = 1;
  ram[32959]  = 1;
  ram[32960]  = 1;
  ram[32961]  = 1;
  ram[32962]  = 1;
  ram[32963]  = 1;
  ram[32964]  = 1;
  ram[32965]  = 1;
  ram[32966]  = 1;
  ram[32967]  = 1;
  ram[32968]  = 1;
  ram[32969]  = 1;
  ram[32970]  = 1;
  ram[32971]  = 1;
  ram[32972]  = 1;
  ram[32973]  = 1;
  ram[32974]  = 1;
  ram[32975]  = 1;
  ram[32976]  = 1;
  ram[32977]  = 1;
  ram[32978]  = 1;
  ram[32979]  = 0;
  ram[32980]  = 1;
  ram[32981]  = 1;
  ram[32982]  = 1;
  ram[32983]  = 1;
  ram[32984]  = 1;
  ram[32985]  = 1;
  ram[32986]  = 1;
  ram[32987]  = 1;
  ram[32988]  = 1;
  ram[32989]  = 1;
  ram[32990]  = 1;
  ram[32991]  = 1;
  ram[32992]  = 1;
  ram[32993]  = 1;
  ram[32994]  = 1;
  ram[32995]  = 1;
  ram[32996]  = 1;
  ram[32997]  = 1;
  ram[32998]  = 1;
  ram[32999]  = 1;
  ram[33000]  = 1;
  ram[33001]  = 1;
  ram[33002]  = 1;
  ram[33003]  = 1;
  ram[33004]  = 1;
  ram[33005]  = 1;
  ram[33006]  = 1;
  ram[33007]  = 1;
  ram[33008]  = 1;
  ram[33009]  = 1;
  ram[33010]  = 1;
  ram[33011]  = 1;
  ram[33012]  = 1;
  ram[33013]  = 1;
  ram[33014]  = 0;
  ram[33015]  = 0;
  ram[33016]  = 1;
  ram[33017]  = 1;
  ram[33018]  = 1;
  ram[33019]  = 0;
  ram[33020]  = 1;
  ram[33021]  = 1;
  ram[33022]  = 1;
  ram[33023]  = 1;
  ram[33024]  = 1;
  ram[33025]  = 1;
  ram[33026]  = 1;
  ram[33027]  = 0;
  ram[33028]  = 1;
  ram[33029]  = 1;
  ram[33030]  = 1;
  ram[33031]  = 1;
  ram[33032]  = 1;
  ram[33033]  = 1;
  ram[33034]  = 1;
  ram[33035]  = 1;
  ram[33036]  = 1;
  ram[33037]  = 1;
  ram[33038]  = 1;
  ram[33039]  = 1;
  ram[33040]  = 1;
  ram[33041]  = 1;
  ram[33042]  = 1;
  ram[33043]  = 1;
  ram[33044]  = 1;
  ram[33045]  = 1;
  ram[33046]  = 1;
  ram[33047]  = 1;
  ram[33048]  = 0;
  ram[33049]  = 1;
  ram[33050]  = 1;
  ram[33051]  = 1;
  ram[33052]  = 1;
  ram[33053]  = 1;
  ram[33054]  = 1;
  ram[33055]  = 1;
  ram[33056]  = 0;
  ram[33057]  = 1;
  ram[33058]  = 1;
  ram[33059]  = 1;
  ram[33060]  = 1;
  ram[33061]  = 1;
  ram[33062]  = 1;
  ram[33063]  = 1;
  ram[33064]  = 1;
  ram[33065]  = 1;
  ram[33066]  = 1;
  ram[33067]  = 1;
  ram[33068]  = 0;
  ram[33069]  = 1;
  ram[33070]  = 1;
  ram[33071]  = 1;
  ram[33072]  = 1;
  ram[33073]  = 1;
  ram[33074]  = 1;
  ram[33075]  = 1;
  ram[33076]  = 1;
  ram[33077]  = 0;
  ram[33078]  = 1;
  ram[33079]  = 1;
  ram[33080]  = 1;
  ram[33081]  = 1;
  ram[33082]  = 1;
  ram[33083]  = 1;
  ram[33084]  = 1;
  ram[33085]  = 1;
  ram[33086]  = 1;
  ram[33087]  = 1;
  ram[33088]  = 0;
  ram[33089]  = 1;
  ram[33090]  = 1;
  ram[33091]  = 1;
  ram[33092]  = 1;
  ram[33093]  = 1;
  ram[33094]  = 0;
  ram[33095]  = 1;
  ram[33096]  = 1;
  ram[33097]  = 1;
  ram[33098]  = 1;
  ram[33099]  = 1;
  ram[33100]  = 1;
  ram[33101]  = 1;
  ram[33102]  = 1;
  ram[33103]  = 1;
  ram[33104]  = 1;
  ram[33105]  = 1;
  ram[33106]  = 1;
  ram[33107]  = 1;
  ram[33108]  = 1;
  ram[33109]  = 1;
  ram[33110]  = 1;
  ram[33111]  = 0;
  ram[33112]  = 1;
  ram[33113]  = 1;
  ram[33114]  = 1;
  ram[33115]  = 1;
  ram[33116]  = 1;
  ram[33117]  = 1;
  ram[33118]  = 1;
  ram[33119]  = 1;
  ram[33120]  = 1;
  ram[33121]  = 1;
  ram[33122]  = 1;
  ram[33123]  = 1;
  ram[33124]  = 0;
  ram[33125]  = 1;
  ram[33126]  = 1;
  ram[33127]  = 1;
  ram[33128]  = 1;
  ram[33129]  = 1;
  ram[33130]  = 0;
  ram[33131]  = 1;
  ram[33132]  = 1;
  ram[33133]  = 1;
  ram[33134]  = 1;
  ram[33135]  = 1;
  ram[33136]  = 1;
  ram[33137]  = 1;
  ram[33138]  = 1;
  ram[33139]  = 1;
  ram[33140]  = 1;
  ram[33141]  = 1;
  ram[33142]  = 1;
  ram[33143]  = 0;
  ram[33144]  = 1;
  ram[33145]  = 1;
  ram[33146]  = 1;
  ram[33147]  = 1;
  ram[33148]  = 1;
  ram[33149]  = 1;
  ram[33150]  = 1;
  ram[33151]  = 1;
  ram[33152]  = 1;
  ram[33153]  = 1;
  ram[33154]  = 1;
  ram[33155]  = 1;
  ram[33156]  = 1;
  ram[33157]  = 1;
  ram[33158]  = 1;
  ram[33159]  = 1;
  ram[33160]  = 1;
  ram[33161]  = 1;
  ram[33162]  = 1;
  ram[33163]  = 1;
  ram[33164]  = 1;
  ram[33165]  = 1;
  ram[33166]  = 1;
  ram[33167]  = 0;
  ram[33168]  = 1;
  ram[33169]  = 1;
  ram[33170]  = 1;
  ram[33171]  = 1;
  ram[33172]  = 1;
  ram[33173]  = 1;
  ram[33174]  = 1;
  ram[33175]  = 1;
  ram[33176]  = 1;
  ram[33177]  = 1;
  ram[33178]  = 1;
  ram[33179]  = 1;
  ram[33180]  = 1;
  ram[33181]  = 1;
  ram[33182]  = 0;
  ram[33183]  = 1;
  ram[33184]  = 1;
  ram[33185]  = 1;
  ram[33186]  = 1;
  ram[33187]  = 1;
  ram[33188]  = 1;
  ram[33189]  = 1;
  ram[33190]  = 1;
  ram[33191]  = 1;
  ram[33192]  = 1;
  ram[33193]  = 0;
  ram[33194]  = 1;
  ram[33195]  = 1;
  ram[33196]  = 1;
  ram[33197]  = 1;
  ram[33198]  = 1;
  ram[33199]  = 1;
  ram[33200]  = 1;
  ram[33201]  = 1;
  ram[33202]  = 1;
  ram[33203]  = 1;
  ram[33204]  = 1;
  ram[33205]  = 0;
  ram[33206]  = 1;
  ram[33207]  = 1;
  ram[33208]  = 1;
  ram[33209]  = 1;
  ram[33210]  = 1;
  ram[33211]  = 0;
  ram[33212]  = 1;
  ram[33213]  = 1;
  ram[33214]  = 0;
  ram[33215]  = 1;
  ram[33216]  = 1;
  ram[33217]  = 1;
  ram[33218]  = 1;
  ram[33219]  = 1;
  ram[33220]  = 1;
  ram[33221]  = 1;
  ram[33222]  = 1;
  ram[33223]  = 1;
  ram[33224]  = 0;
  ram[33225]  = 1;
  ram[33226]  = 1;
  ram[33227]  = 1;
  ram[33228]  = 1;
  ram[33229]  = 1;
  ram[33230]  = 1;
  ram[33231]  = 1;
  ram[33232]  = 1;
  ram[33233]  = 1;
  ram[33234]  = 1;
  ram[33235]  = 0;
  ram[33236]  = 0;
  ram[33237]  = 1;
  ram[33238]  = 1;
  ram[33239]  = 0;
  ram[33240]  = 1;
  ram[33241]  = 1;
  ram[33242]  = 1;
  ram[33243]  = 1;
  ram[33244]  = 1;
  ram[33245]  = 1;
  ram[33246]  = 1;
  ram[33247]  = 1;
  ram[33248]  = 1;
  ram[33249]  = 1;
  ram[33250]  = 1;
  ram[33251]  = 1;
  ram[33252]  = 1;
  ram[33253]  = 1;
  ram[33254]  = 1;
  ram[33255]  = 1;
  ram[33256]  = 1;
  ram[33257]  = 1;
  ram[33258]  = 1;
  ram[33259]  = 0;
  ram[33260]  = 1;
  ram[33261]  = 1;
  ram[33262]  = 1;
  ram[33263]  = 1;
  ram[33264]  = 1;
  ram[33265]  = 1;
  ram[33266]  = 1;
  ram[33267]  = 1;
  ram[33268]  = 1;
  ram[33269]  = 1;
  ram[33270]  = 1;
  ram[33271]  = 1;
  ram[33272]  = 1;
  ram[33273]  = 1;
  ram[33274]  = 1;
  ram[33275]  = 0;
  ram[33276]  = 1;
  ram[33277]  = 1;
  ram[33278]  = 1;
  ram[33279]  = 0;
  ram[33280]  = 1;
  ram[33281]  = 1;
  ram[33282]  = 1;
  ram[33283]  = 1;
  ram[33284]  = 1;
  ram[33285]  = 1;
  ram[33286]  = 1;
  ram[33287]  = 1;
  ram[33288]  = 1;
  ram[33289]  = 1;
  ram[33290]  = 1;
  ram[33291]  = 1;
  ram[33292]  = 1;
  ram[33293]  = 1;
  ram[33294]  = 1;
  ram[33295]  = 1;
  ram[33296]  = 1;
  ram[33297]  = 1;
  ram[33298]  = 1;
  ram[33299]  = 1;
  ram[33300]  = 1;
  ram[33301]  = 1;
  ram[33302]  = 1;
  ram[33303]  = 1;
  ram[33304]  = 1;
  ram[33305]  = 1;
  ram[33306]  = 1;
  ram[33307]  = 1;
  ram[33308]  = 1;
  ram[33309]  = 1;
  ram[33310]  = 1;
  ram[33311]  = 1;
  ram[33312]  = 1;
  ram[33313]  = 1;
  ram[33314]  = 1;
  ram[33315]  = 0;
  ram[33316]  = 1;
  ram[33317]  = 1;
  ram[33318]  = 1;
  ram[33319]  = 0;
  ram[33320]  = 1;
  ram[33321]  = 1;
  ram[33322]  = 1;
  ram[33323]  = 1;
  ram[33324]  = 1;
  ram[33325]  = 0;
  ram[33326]  = 0;
  ram[33327]  = 0;
  ram[33328]  = 0;
  ram[33329]  = 0;
  ram[33330]  = 1;
  ram[33331]  = 1;
  ram[33332]  = 1;
  ram[33333]  = 1;
  ram[33334]  = 0;
  ram[33335]  = 0;
  ram[33336]  = 1;
  ram[33337]  = 1;
  ram[33338]  = 1;
  ram[33339]  = 1;
  ram[33340]  = 1;
  ram[33341]  = 0;
  ram[33342]  = 1;
  ram[33343]  = 1;
  ram[33344]  = 1;
  ram[33345]  = 0;
  ram[33346]  = 1;
  ram[33347]  = 0;
  ram[33348]  = 0;
  ram[33349]  = 1;
  ram[33350]  = 1;
  ram[33351]  = 1;
  ram[33352]  = 1;
  ram[33353]  = 1;
  ram[33354]  = 1;
  ram[33355]  = 1;
  ram[33356]  = 0;
  ram[33357]  = 1;
  ram[33358]  = 1;
  ram[33359]  = 1;
  ram[33360]  = 1;
  ram[33361]  = 1;
  ram[33362]  = 1;
  ram[33363]  = 1;
  ram[33364]  = 1;
  ram[33365]  = 1;
  ram[33366]  = 1;
  ram[33367]  = 0;
  ram[33368]  = 0;
  ram[33369]  = 0;
  ram[33370]  = 0;
  ram[33371]  = 1;
  ram[33372]  = 1;
  ram[33373]  = 1;
  ram[33374]  = 1;
  ram[33375]  = 0;
  ram[33376]  = 0;
  ram[33377]  = 0;
  ram[33378]  = 0;
  ram[33379]  = 0;
  ram[33380]  = 1;
  ram[33381]  = 1;
  ram[33382]  = 1;
  ram[33383]  = 1;
  ram[33384]  = 1;
  ram[33385]  = 0;
  ram[33386]  = 1;
  ram[33387]  = 0;
  ram[33388]  = 0;
  ram[33389]  = 1;
  ram[33390]  = 1;
  ram[33391]  = 1;
  ram[33392]  = 0;
  ram[33393]  = 0;
  ram[33394]  = 0;
  ram[33395]  = 0;
  ram[33396]  = 0;
  ram[33397]  = 1;
  ram[33398]  = 1;
  ram[33399]  = 1;
  ram[33400]  = 1;
  ram[33401]  = 1;
  ram[33402]  = 1;
  ram[33403]  = 1;
  ram[33404]  = 1;
  ram[33405]  = 0;
  ram[33406]  = 0;
  ram[33407]  = 1;
  ram[33408]  = 1;
  ram[33409]  = 1;
  ram[33410]  = 0;
  ram[33411]  = 0;
  ram[33412]  = 0;
  ram[33413]  = 0;
  ram[33414]  = 1;
  ram[33415]  = 1;
  ram[33416]  = 1;
  ram[33417]  = 1;
  ram[33418]  = 1;
  ram[33419]  = 1;
  ram[33420]  = 1;
  ram[33421]  = 1;
  ram[33422]  = 0;
  ram[33423]  = 0;
  ram[33424]  = 0;
  ram[33425]  = 0;
  ram[33426]  = 0;
  ram[33427]  = 1;
  ram[33428]  = 1;
  ram[33429]  = 1;
  ram[33430]  = 0;
  ram[33431]  = 1;
  ram[33432]  = 0;
  ram[33433]  = 0;
  ram[33434]  = 0;
  ram[33435]  = 0;
  ram[33436]  = 1;
  ram[33437]  = 1;
  ram[33438]  = 1;
  ram[33439]  = 1;
  ram[33440]  = 1;
  ram[33441]  = 0;
  ram[33442]  = 0;
  ram[33443]  = 0;
  ram[33444]  = 0;
  ram[33445]  = 0;
  ram[33446]  = 1;
  ram[33447]  = 1;
  ram[33448]  = 1;
  ram[33449]  = 0;
  ram[33450]  = 0;
  ram[33451]  = 1;
  ram[33452]  = 1;
  ram[33453]  = 1;
  ram[33454]  = 1;
  ram[33455]  = 0;
  ram[33456]  = 1;
  ram[33457]  = 1;
  ram[33458]  = 1;
  ram[33459]  = 1;
  ram[33460]  = 1;
  ram[33461]  = 0;
  ram[33462]  = 1;
  ram[33463]  = 1;
  ram[33464]  = 0;
  ram[33465]  = 1;
  ram[33466]  = 0;
  ram[33467]  = 0;
  ram[33468]  = 0;
  ram[33469]  = 0;
  ram[33470]  = 1;
  ram[33471]  = 1;
  ram[33472]  = 1;
  ram[33473]  = 1;
  ram[33474]  = 1;
  ram[33475]  = 1;
  ram[33476]  = 1;
  ram[33477]  = 1;
  ram[33478]  = 1;
  ram[33479]  = 1;
  ram[33480]  = 0;
  ram[33481]  = 0;
  ram[33482]  = 0;
  ram[33483]  = 0;
  ram[33484]  = 0;
  ram[33485]  = 1;
  ram[33486]  = 1;
  ram[33487]  = 1;
  ram[33488]  = 1;
  ram[33489]  = 0;
  ram[33490]  = 0;
  ram[33491]  = 1;
  ram[33492]  = 0;
  ram[33493]  = 0;
  ram[33494]  = 0;
  ram[33495]  = 0;
  ram[33496]  = 1;
  ram[33497]  = 1;
  ram[33498]  = 1;
  ram[33499]  = 1;
  ram[33500]  = 1;
  ram[33501]  = 1;
  ram[33502]  = 1;
  ram[33503]  = 1;
  ram[33504]  = 0;
  ram[33505]  = 0;
  ram[33506]  = 0;
  ram[33507]  = 0;
  ram[33508]  = 0;
  ram[33509]  = 1;
  ram[33510]  = 1;
  ram[33511]  = 0;
  ram[33512]  = 1;
  ram[33513]  = 0;
  ram[33514]  = 0;
  ram[33515]  = 0;
  ram[33516]  = 0;
  ram[33517]  = 1;
  ram[33518]  = 1;
  ram[33519]  = 1;
  ram[33520]  = 1;
  ram[33521]  = 1;
  ram[33522]  = 0;
  ram[33523]  = 0;
  ram[33524]  = 0;
  ram[33525]  = 0;
  ram[33526]  = 0;
  ram[33527]  = 1;
  ram[33528]  = 1;
  ram[33529]  = 1;
  ram[33530]  = 1;
  ram[33531]  = 1;
  ram[33532]  = 1;
  ram[33533]  = 1;
  ram[33534]  = 1;
  ram[33535]  = 0;
  ram[33536]  = 0;
  ram[33537]  = 1;
  ram[33538]  = 0;
  ram[33539]  = 0;
  ram[33540]  = 0;
  ram[33541]  = 0;
  ram[33542]  = 1;
  ram[33543]  = 1;
  ram[33544]  = 1;
  ram[33545]  = 1;
  ram[33546]  = 1;
  ram[33547]  = 1;
  ram[33548]  = 0;
  ram[33549]  = 0;
  ram[33550]  = 0;
  ram[33551]  = 0;
  ram[33552]  = 1;
  ram[33553]  = 1;
  ram[33554]  = 1;
  ram[33555]  = 1;
  ram[33556]  = 1;
  ram[33557]  = 0;
  ram[33558]  = 0;
  ram[33559]  = 0;
  ram[33560]  = 0;
  ram[33561]  = 0;
  ram[33562]  = 1;
  ram[33563]  = 1;
  ram[33564]  = 1;
  ram[33565]  = 1;
  ram[33566]  = 0;
  ram[33567]  = 1;
  ram[33568]  = 0;
  ram[33569]  = 0;
  ram[33570]  = 0;
  ram[33571]  = 1;
  ram[33572]  = 1;
  ram[33573]  = 1;
  ram[33574]  = 0;
  ram[33575]  = 0;
  ram[33576]  = 0;
  ram[33577]  = 0;
  ram[33578]  = 1;
  ram[33579]  = 0;
  ram[33580]  = 1;
  ram[33581]  = 1;
  ram[33582]  = 1;
  ram[33583]  = 1;
  ram[33584]  = 1;
  ram[33585]  = 1;
  ram[33586]  = 1;
  ram[33587]  = 1;
  ram[33588]  = 1;
  ram[33589]  = 1;
  ram[33590]  = 1;
  ram[33591]  = 1;
  ram[33592]  = 1;
  ram[33593]  = 1;
  ram[33594]  = 1;
  ram[33595]  = 1;
  ram[33596]  = 1;
  ram[33597]  = 1;
  ram[33598]  = 1;
  ram[33599]  = 1;
  ram[33600]  = 1;
  ram[33601]  = 1;
  ram[33602]  = 1;
  ram[33603]  = 1;
  ram[33604]  = 1;
  ram[33605]  = 1;
  ram[33606]  = 1;
  ram[33607]  = 1;
  ram[33608]  = 1;
  ram[33609]  = 1;
  ram[33610]  = 1;
  ram[33611]  = 1;
  ram[33612]  = 1;
  ram[33613]  = 1;
  ram[33614]  = 1;
  ram[33615]  = 0;
  ram[33616]  = 1;
  ram[33617]  = 1;
  ram[33618]  = 0;
  ram[33619]  = 0;
  ram[33620]  = 1;
  ram[33621]  = 1;
  ram[33622]  = 1;
  ram[33623]  = 1;
  ram[33624]  = 1;
  ram[33625]  = 0;
  ram[33626]  = 0;
  ram[33627]  = 1;
  ram[33628]  = 1;
  ram[33629]  = 0;
  ram[33630]  = 0;
  ram[33631]  = 1;
  ram[33632]  = 1;
  ram[33633]  = 1;
  ram[33634]  = 0;
  ram[33635]  = 0;
  ram[33636]  = 1;
  ram[33637]  = 1;
  ram[33638]  = 1;
  ram[33639]  = 1;
  ram[33640]  = 1;
  ram[33641]  = 0;
  ram[33642]  = 1;
  ram[33643]  = 1;
  ram[33644]  = 1;
  ram[33645]  = 0;
  ram[33646]  = 0;
  ram[33647]  = 0;
  ram[33648]  = 1;
  ram[33649]  = 1;
  ram[33650]  = 1;
  ram[33651]  = 1;
  ram[33652]  = 1;
  ram[33653]  = 1;
  ram[33654]  = 1;
  ram[33655]  = 1;
  ram[33656]  = 0;
  ram[33657]  = 1;
  ram[33658]  = 1;
  ram[33659]  = 1;
  ram[33660]  = 1;
  ram[33661]  = 1;
  ram[33662]  = 1;
  ram[33663]  = 1;
  ram[33664]  = 1;
  ram[33665]  = 1;
  ram[33666]  = 0;
  ram[33667]  = 0;
  ram[33668]  = 1;
  ram[33669]  = 1;
  ram[33670]  = 0;
  ram[33671]  = 0;
  ram[33672]  = 1;
  ram[33673]  = 1;
  ram[33674]  = 1;
  ram[33675]  = 0;
  ram[33676]  = 0;
  ram[33677]  = 1;
  ram[33678]  = 1;
  ram[33679]  = 0;
  ram[33680]  = 0;
  ram[33681]  = 1;
  ram[33682]  = 1;
  ram[33683]  = 1;
  ram[33684]  = 1;
  ram[33685]  = 0;
  ram[33686]  = 0;
  ram[33687]  = 1;
  ram[33688]  = 1;
  ram[33689]  = 1;
  ram[33690]  = 1;
  ram[33691]  = 0;
  ram[33692]  = 0;
  ram[33693]  = 1;
  ram[33694]  = 1;
  ram[33695]  = 0;
  ram[33696]  = 0;
  ram[33697]  = 1;
  ram[33698]  = 1;
  ram[33699]  = 1;
  ram[33700]  = 1;
  ram[33701]  = 1;
  ram[33702]  = 1;
  ram[33703]  = 1;
  ram[33704]  = 1;
  ram[33705]  = 0;
  ram[33706]  = 0;
  ram[33707]  = 1;
  ram[33708]  = 1;
  ram[33709]  = 0;
  ram[33710]  = 0;
  ram[33711]  = 1;
  ram[33712]  = 1;
  ram[33713]  = 0;
  ram[33714]  = 0;
  ram[33715]  = 1;
  ram[33716]  = 1;
  ram[33717]  = 1;
  ram[33718]  = 1;
  ram[33719]  = 1;
  ram[33720]  = 1;
  ram[33721]  = 1;
  ram[33722]  = 0;
  ram[33723]  = 1;
  ram[33724]  = 1;
  ram[33725]  = 1;
  ram[33726]  = 0;
  ram[33727]  = 1;
  ram[33728]  = 1;
  ram[33729]  = 1;
  ram[33730]  = 0;
  ram[33731]  = 0;
  ram[33732]  = 0;
  ram[33733]  = 1;
  ram[33734]  = 1;
  ram[33735]  = 0;
  ram[33736]  = 0;
  ram[33737]  = 1;
  ram[33738]  = 1;
  ram[33739]  = 1;
  ram[33740]  = 1;
  ram[33741]  = 0;
  ram[33742]  = 0;
  ram[33743]  = 1;
  ram[33744]  = 1;
  ram[33745]  = 0;
  ram[33746]  = 0;
  ram[33747]  = 1;
  ram[33748]  = 1;
  ram[33749]  = 1;
  ram[33750]  = 0;
  ram[33751]  = 1;
  ram[33752]  = 1;
  ram[33753]  = 1;
  ram[33754]  = 1;
  ram[33755]  = 0;
  ram[33756]  = 1;
  ram[33757]  = 1;
  ram[33758]  = 1;
  ram[33759]  = 1;
  ram[33760]  = 0;
  ram[33761]  = 0;
  ram[33762]  = 1;
  ram[33763]  = 1;
  ram[33764]  = 0;
  ram[33765]  = 0;
  ram[33766]  = 0;
  ram[33767]  = 1;
  ram[33768]  = 1;
  ram[33769]  = 0;
  ram[33770]  = 1;
  ram[33771]  = 1;
  ram[33772]  = 1;
  ram[33773]  = 1;
  ram[33774]  = 1;
  ram[33775]  = 1;
  ram[33776]  = 1;
  ram[33777]  = 1;
  ram[33778]  = 1;
  ram[33779]  = 1;
  ram[33780]  = 0;
  ram[33781]  = 0;
  ram[33782]  = 1;
  ram[33783]  = 1;
  ram[33784]  = 0;
  ram[33785]  = 0;
  ram[33786]  = 1;
  ram[33787]  = 1;
  ram[33788]  = 1;
  ram[33789]  = 1;
  ram[33790]  = 0;
  ram[33791]  = 0;
  ram[33792]  = 1;
  ram[33793]  = 1;
  ram[33794]  = 0;
  ram[33795]  = 0;
  ram[33796]  = 1;
  ram[33797]  = 1;
  ram[33798]  = 1;
  ram[33799]  = 1;
  ram[33800]  = 1;
  ram[33801]  = 1;
  ram[33802]  = 1;
  ram[33803]  = 1;
  ram[33804]  = 1;
  ram[33805]  = 0;
  ram[33806]  = 0;
  ram[33807]  = 0;
  ram[33808]  = 1;
  ram[33809]  = 1;
  ram[33810]  = 1;
  ram[33811]  = 0;
  ram[33812]  = 0;
  ram[33813]  = 0;
  ram[33814]  = 1;
  ram[33815]  = 0;
  ram[33816]  = 0;
  ram[33817]  = 1;
  ram[33818]  = 1;
  ram[33819]  = 1;
  ram[33820]  = 1;
  ram[33821]  = 0;
  ram[33822]  = 0;
  ram[33823]  = 1;
  ram[33824]  = 1;
  ram[33825]  = 0;
  ram[33826]  = 0;
  ram[33827]  = 1;
  ram[33828]  = 1;
  ram[33829]  = 1;
  ram[33830]  = 1;
  ram[33831]  = 1;
  ram[33832]  = 1;
  ram[33833]  = 1;
  ram[33834]  = 1;
  ram[33835]  = 0;
  ram[33836]  = 0;
  ram[33837]  = 0;
  ram[33838]  = 0;
  ram[33839]  = 1;
  ram[33840]  = 1;
  ram[33841]  = 0;
  ram[33842]  = 0;
  ram[33843]  = 1;
  ram[33844]  = 1;
  ram[33845]  = 1;
  ram[33846]  = 1;
  ram[33847]  = 0;
  ram[33848]  = 0;
  ram[33849]  = 1;
  ram[33850]  = 1;
  ram[33851]  = 0;
  ram[33852]  = 0;
  ram[33853]  = 1;
  ram[33854]  = 1;
  ram[33855]  = 1;
  ram[33856]  = 1;
  ram[33857]  = 0;
  ram[33858]  = 0;
  ram[33859]  = 1;
  ram[33860]  = 1;
  ram[33861]  = 0;
  ram[33862]  = 0;
  ram[33863]  = 1;
  ram[33864]  = 1;
  ram[33865]  = 1;
  ram[33866]  = 0;
  ram[33867]  = 1;
  ram[33868]  = 0;
  ram[33869]  = 1;
  ram[33870]  = 1;
  ram[33871]  = 1;
  ram[33872]  = 1;
  ram[33873]  = 0;
  ram[33874]  = 0;
  ram[33875]  = 1;
  ram[33876]  = 1;
  ram[33877]  = 0;
  ram[33878]  = 0;
  ram[33879]  = 0;
  ram[33880]  = 1;
  ram[33881]  = 1;
  ram[33882]  = 1;
  ram[33883]  = 1;
  ram[33884]  = 1;
  ram[33885]  = 1;
  ram[33886]  = 1;
  ram[33887]  = 1;
  ram[33888]  = 1;
  ram[33889]  = 1;
  ram[33890]  = 1;
  ram[33891]  = 1;
  ram[33892]  = 1;
  ram[33893]  = 1;
  ram[33894]  = 1;
  ram[33895]  = 1;
  ram[33896]  = 1;
  ram[33897]  = 1;
  ram[33898]  = 1;
  ram[33899]  = 1;
  ram[33900]  = 1;
  ram[33901]  = 1;
  ram[33902]  = 1;
  ram[33903]  = 1;
  ram[33904]  = 1;
  ram[33905]  = 1;
  ram[33906]  = 1;
  ram[33907]  = 1;
  ram[33908]  = 1;
  ram[33909]  = 1;
  ram[33910]  = 1;
  ram[33911]  = 1;
  ram[33912]  = 1;
  ram[33913]  = 1;
  ram[33914]  = 1;
  ram[33915]  = 0;
  ram[33916]  = 0;
  ram[33917]  = 1;
  ram[33918]  = 0;
  ram[33919]  = 1;
  ram[33920]  = 1;
  ram[33921]  = 1;
  ram[33922]  = 1;
  ram[33923]  = 1;
  ram[33924]  = 0;
  ram[33925]  = 0;
  ram[33926]  = 1;
  ram[33927]  = 1;
  ram[33928]  = 1;
  ram[33929]  = 1;
  ram[33930]  = 0;
  ram[33931]  = 1;
  ram[33932]  = 1;
  ram[33933]  = 1;
  ram[33934]  = 0;
  ram[33935]  = 0;
  ram[33936]  = 1;
  ram[33937]  = 1;
  ram[33938]  = 1;
  ram[33939]  = 1;
  ram[33940]  = 1;
  ram[33941]  = 0;
  ram[33942]  = 1;
  ram[33943]  = 1;
  ram[33944]  = 1;
  ram[33945]  = 0;
  ram[33946]  = 0;
  ram[33947]  = 1;
  ram[33948]  = 1;
  ram[33949]  = 1;
  ram[33950]  = 1;
  ram[33951]  = 1;
  ram[33952]  = 1;
  ram[33953]  = 1;
  ram[33954]  = 1;
  ram[33955]  = 1;
  ram[33956]  = 0;
  ram[33957]  = 0;
  ram[33958]  = 1;
  ram[33959]  = 1;
  ram[33960]  = 1;
  ram[33961]  = 1;
  ram[33962]  = 1;
  ram[33963]  = 1;
  ram[33964]  = 1;
  ram[33965]  = 1;
  ram[33966]  = 0;
  ram[33967]  = 1;
  ram[33968]  = 1;
  ram[33969]  = 1;
  ram[33970]  = 1;
  ram[33971]  = 0;
  ram[33972]  = 1;
  ram[33973]  = 1;
  ram[33974]  = 0;
  ram[33975]  = 0;
  ram[33976]  = 1;
  ram[33977]  = 1;
  ram[33978]  = 1;
  ram[33979]  = 1;
  ram[33980]  = 0;
  ram[33981]  = 0;
  ram[33982]  = 1;
  ram[33983]  = 1;
  ram[33984]  = 1;
  ram[33985]  = 0;
  ram[33986]  = 0;
  ram[33987]  = 1;
  ram[33988]  = 1;
  ram[33989]  = 1;
  ram[33990]  = 1;
  ram[33991]  = 0;
  ram[33992]  = 1;
  ram[33993]  = 1;
  ram[33994]  = 1;
  ram[33995]  = 1;
  ram[33996]  = 0;
  ram[33997]  = 0;
  ram[33998]  = 1;
  ram[33999]  = 1;
  ram[34000]  = 1;
  ram[34001]  = 1;
  ram[34002]  = 1;
  ram[34003]  = 1;
  ram[34004]  = 1;
  ram[34005]  = 0;
  ram[34006]  = 0;
  ram[34007]  = 1;
  ram[34008]  = 1;
  ram[34009]  = 0;
  ram[34010]  = 1;
  ram[34011]  = 1;
  ram[34012]  = 1;
  ram[34013]  = 1;
  ram[34014]  = 0;
  ram[34015]  = 1;
  ram[34016]  = 1;
  ram[34017]  = 1;
  ram[34018]  = 1;
  ram[34019]  = 1;
  ram[34020]  = 1;
  ram[34021]  = 1;
  ram[34022]  = 0;
  ram[34023]  = 1;
  ram[34024]  = 1;
  ram[34025]  = 1;
  ram[34026]  = 0;
  ram[34027]  = 0;
  ram[34028]  = 1;
  ram[34029]  = 1;
  ram[34030]  = 0;
  ram[34031]  = 0;
  ram[34032]  = 1;
  ram[34033]  = 1;
  ram[34034]  = 1;
  ram[34035]  = 0;
  ram[34036]  = 0;
  ram[34037]  = 1;
  ram[34038]  = 1;
  ram[34039]  = 1;
  ram[34040]  = 0;
  ram[34041]  = 0;
  ram[34042]  = 1;
  ram[34043]  = 1;
  ram[34044]  = 1;
  ram[34045]  = 1;
  ram[34046]  = 0;
  ram[34047]  = 0;
  ram[34048]  = 1;
  ram[34049]  = 1;
  ram[34050]  = 0;
  ram[34051]  = 1;
  ram[34052]  = 1;
  ram[34053]  = 1;
  ram[34054]  = 1;
  ram[34055]  = 0;
  ram[34056]  = 0;
  ram[34057]  = 1;
  ram[34058]  = 1;
  ram[34059]  = 1;
  ram[34060]  = 0;
  ram[34061]  = 1;
  ram[34062]  = 1;
  ram[34063]  = 1;
  ram[34064]  = 0;
  ram[34065]  = 0;
  ram[34066]  = 1;
  ram[34067]  = 1;
  ram[34068]  = 1;
  ram[34069]  = 0;
  ram[34070]  = 0;
  ram[34071]  = 1;
  ram[34072]  = 1;
  ram[34073]  = 1;
  ram[34074]  = 1;
  ram[34075]  = 1;
  ram[34076]  = 1;
  ram[34077]  = 1;
  ram[34078]  = 1;
  ram[34079]  = 0;
  ram[34080]  = 0;
  ram[34081]  = 1;
  ram[34082]  = 1;
  ram[34083]  = 1;
  ram[34084]  = 1;
  ram[34085]  = 0;
  ram[34086]  = 1;
  ram[34087]  = 1;
  ram[34088]  = 1;
  ram[34089]  = 1;
  ram[34090]  = 0;
  ram[34091]  = 0;
  ram[34092]  = 1;
  ram[34093]  = 1;
  ram[34094]  = 1;
  ram[34095]  = 0;
  ram[34096]  = 0;
  ram[34097]  = 1;
  ram[34098]  = 1;
  ram[34099]  = 1;
  ram[34100]  = 1;
  ram[34101]  = 1;
  ram[34102]  = 1;
  ram[34103]  = 1;
  ram[34104]  = 1;
  ram[34105]  = 0;
  ram[34106]  = 1;
  ram[34107]  = 1;
  ram[34108]  = 1;
  ram[34109]  = 1;
  ram[34110]  = 1;
  ram[34111]  = 0;
  ram[34112]  = 0;
  ram[34113]  = 1;
  ram[34114]  = 1;
  ram[34115]  = 1;
  ram[34116]  = 0;
  ram[34117]  = 0;
  ram[34118]  = 1;
  ram[34119]  = 1;
  ram[34120]  = 1;
  ram[34121]  = 0;
  ram[34122]  = 1;
  ram[34123]  = 1;
  ram[34124]  = 1;
  ram[34125]  = 1;
  ram[34126]  = 0;
  ram[34127]  = 0;
  ram[34128]  = 1;
  ram[34129]  = 1;
  ram[34130]  = 1;
  ram[34131]  = 1;
  ram[34132]  = 1;
  ram[34133]  = 1;
  ram[34134]  = 1;
  ram[34135]  = 0;
  ram[34136]  = 0;
  ram[34137]  = 0;
  ram[34138]  = 1;
  ram[34139]  = 1;
  ram[34140]  = 1;
  ram[34141]  = 1;
  ram[34142]  = 0;
  ram[34143]  = 1;
  ram[34144]  = 1;
  ram[34145]  = 1;
  ram[34146]  = 0;
  ram[34147]  = 0;
  ram[34148]  = 1;
  ram[34149]  = 1;
  ram[34150]  = 1;
  ram[34151]  = 1;
  ram[34152]  = 0;
  ram[34153]  = 0;
  ram[34154]  = 1;
  ram[34155]  = 1;
  ram[34156]  = 1;
  ram[34157]  = 0;
  ram[34158]  = 1;
  ram[34159]  = 1;
  ram[34160]  = 1;
  ram[34161]  = 0;
  ram[34162]  = 0;
  ram[34163]  = 1;
  ram[34164]  = 1;
  ram[34165]  = 1;
  ram[34166]  = 0;
  ram[34167]  = 0;
  ram[34168]  = 1;
  ram[34169]  = 1;
  ram[34170]  = 1;
  ram[34171]  = 1;
  ram[34172]  = 1;
  ram[34173]  = 0;
  ram[34174]  = 1;
  ram[34175]  = 1;
  ram[34176]  = 1;
  ram[34177]  = 1;
  ram[34178]  = 0;
  ram[34179]  = 0;
  ram[34180]  = 1;
  ram[34181]  = 1;
  ram[34182]  = 1;
  ram[34183]  = 1;
  ram[34184]  = 1;
  ram[34185]  = 1;
  ram[34186]  = 1;
  ram[34187]  = 1;
  ram[34188]  = 1;
  ram[34189]  = 1;
  ram[34190]  = 1;
  ram[34191]  = 1;
  ram[34192]  = 1;
  ram[34193]  = 1;
  ram[34194]  = 1;
  ram[34195]  = 1;
  ram[34196]  = 1;
  ram[34197]  = 1;
  ram[34198]  = 1;
  ram[34199]  = 1;
  ram[34200]  = 1;
  ram[34201]  = 1;
  ram[34202]  = 1;
  ram[34203]  = 1;
  ram[34204]  = 1;
  ram[34205]  = 1;
  ram[34206]  = 1;
  ram[34207]  = 1;
  ram[34208]  = 1;
  ram[34209]  = 1;
  ram[34210]  = 1;
  ram[34211]  = 1;
  ram[34212]  = 1;
  ram[34213]  = 1;
  ram[34214]  = 1;
  ram[34215]  = 1;
  ram[34216]  = 0;
  ram[34217]  = 1;
  ram[34218]  = 0;
  ram[34219]  = 1;
  ram[34220]  = 1;
  ram[34221]  = 1;
  ram[34222]  = 1;
  ram[34223]  = 1;
  ram[34224]  = 0;
  ram[34225]  = 1;
  ram[34226]  = 1;
  ram[34227]  = 1;
  ram[34228]  = 1;
  ram[34229]  = 1;
  ram[34230]  = 0;
  ram[34231]  = 0;
  ram[34232]  = 1;
  ram[34233]  = 1;
  ram[34234]  = 0;
  ram[34235]  = 0;
  ram[34236]  = 1;
  ram[34237]  = 1;
  ram[34238]  = 1;
  ram[34239]  = 1;
  ram[34240]  = 1;
  ram[34241]  = 0;
  ram[34242]  = 1;
  ram[34243]  = 1;
  ram[34244]  = 1;
  ram[34245]  = 0;
  ram[34246]  = 1;
  ram[34247]  = 1;
  ram[34248]  = 1;
  ram[34249]  = 1;
  ram[34250]  = 1;
  ram[34251]  = 1;
  ram[34252]  = 1;
  ram[34253]  = 1;
  ram[34254]  = 1;
  ram[34255]  = 1;
  ram[34256]  = 1;
  ram[34257]  = 0;
  ram[34258]  = 0;
  ram[34259]  = 1;
  ram[34260]  = 1;
  ram[34261]  = 1;
  ram[34262]  = 1;
  ram[34263]  = 1;
  ram[34264]  = 1;
  ram[34265]  = 0;
  ram[34266]  = 0;
  ram[34267]  = 1;
  ram[34268]  = 1;
  ram[34269]  = 1;
  ram[34270]  = 1;
  ram[34271]  = 0;
  ram[34272]  = 1;
  ram[34273]  = 1;
  ram[34274]  = 0;
  ram[34275]  = 1;
  ram[34276]  = 1;
  ram[34277]  = 1;
  ram[34278]  = 1;
  ram[34279]  = 1;
  ram[34280]  = 1;
  ram[34281]  = 0;
  ram[34282]  = 1;
  ram[34283]  = 1;
  ram[34284]  = 1;
  ram[34285]  = 0;
  ram[34286]  = 1;
  ram[34287]  = 1;
  ram[34288]  = 1;
  ram[34289]  = 1;
  ram[34290]  = 1;
  ram[34291]  = 0;
  ram[34292]  = 1;
  ram[34293]  = 1;
  ram[34294]  = 1;
  ram[34295]  = 1;
  ram[34296]  = 1;
  ram[34297]  = 0;
  ram[34298]  = 1;
  ram[34299]  = 1;
  ram[34300]  = 1;
  ram[34301]  = 1;
  ram[34302]  = 1;
  ram[34303]  = 1;
  ram[34304]  = 1;
  ram[34305]  = 0;
  ram[34306]  = 0;
  ram[34307]  = 1;
  ram[34308]  = 1;
  ram[34309]  = 0;
  ram[34310]  = 1;
  ram[34311]  = 1;
  ram[34312]  = 1;
  ram[34313]  = 1;
  ram[34314]  = 1;
  ram[34315]  = 1;
  ram[34316]  = 1;
  ram[34317]  = 1;
  ram[34318]  = 1;
  ram[34319]  = 1;
  ram[34320]  = 1;
  ram[34321]  = 1;
  ram[34322]  = 0;
  ram[34323]  = 1;
  ram[34324]  = 1;
  ram[34325]  = 1;
  ram[34326]  = 1;
  ram[34327]  = 1;
  ram[34328]  = 1;
  ram[34329]  = 1;
  ram[34330]  = 0;
  ram[34331]  = 1;
  ram[34332]  = 1;
  ram[34333]  = 1;
  ram[34334]  = 1;
  ram[34335]  = 1;
  ram[34336]  = 0;
  ram[34337]  = 1;
  ram[34338]  = 1;
  ram[34339]  = 1;
  ram[34340]  = 0;
  ram[34341]  = 1;
  ram[34342]  = 1;
  ram[34343]  = 1;
  ram[34344]  = 1;
  ram[34345]  = 1;
  ram[34346]  = 0;
  ram[34347]  = 0;
  ram[34348]  = 1;
  ram[34349]  = 1;
  ram[34350]  = 0;
  ram[34351]  = 1;
  ram[34352]  = 1;
  ram[34353]  = 1;
  ram[34354]  = 0;
  ram[34355]  = 0;
  ram[34356]  = 0;
  ram[34357]  = 1;
  ram[34358]  = 1;
  ram[34359]  = 1;
  ram[34360]  = 0;
  ram[34361]  = 1;
  ram[34362]  = 1;
  ram[34363]  = 1;
  ram[34364]  = 0;
  ram[34365]  = 1;
  ram[34366]  = 1;
  ram[34367]  = 1;
  ram[34368]  = 1;
  ram[34369]  = 1;
  ram[34370]  = 0;
  ram[34371]  = 1;
  ram[34372]  = 1;
  ram[34373]  = 1;
  ram[34374]  = 1;
  ram[34375]  = 1;
  ram[34376]  = 1;
  ram[34377]  = 1;
  ram[34378]  = 1;
  ram[34379]  = 0;
  ram[34380]  = 1;
  ram[34381]  = 1;
  ram[34382]  = 1;
  ram[34383]  = 1;
  ram[34384]  = 1;
  ram[34385]  = 0;
  ram[34386]  = 0;
  ram[34387]  = 1;
  ram[34388]  = 1;
  ram[34389]  = 1;
  ram[34390]  = 0;
  ram[34391]  = 1;
  ram[34392]  = 1;
  ram[34393]  = 1;
  ram[34394]  = 1;
  ram[34395]  = 0;
  ram[34396]  = 0;
  ram[34397]  = 1;
  ram[34398]  = 1;
  ram[34399]  = 1;
  ram[34400]  = 1;
  ram[34401]  = 1;
  ram[34402]  = 1;
  ram[34403]  = 1;
  ram[34404]  = 1;
  ram[34405]  = 0;
  ram[34406]  = 1;
  ram[34407]  = 1;
  ram[34408]  = 1;
  ram[34409]  = 1;
  ram[34410]  = 1;
  ram[34411]  = 0;
  ram[34412]  = 1;
  ram[34413]  = 1;
  ram[34414]  = 1;
  ram[34415]  = 1;
  ram[34416]  = 1;
  ram[34417]  = 0;
  ram[34418]  = 1;
  ram[34419]  = 1;
  ram[34420]  = 1;
  ram[34421]  = 0;
  ram[34422]  = 1;
  ram[34423]  = 1;
  ram[34424]  = 1;
  ram[34425]  = 1;
  ram[34426]  = 1;
  ram[34427]  = 0;
  ram[34428]  = 1;
  ram[34429]  = 1;
  ram[34430]  = 1;
  ram[34431]  = 1;
  ram[34432]  = 1;
  ram[34433]  = 1;
  ram[34434]  = 1;
  ram[34435]  = 1;
  ram[34436]  = 0;
  ram[34437]  = 1;
  ram[34438]  = 1;
  ram[34439]  = 1;
  ram[34440]  = 1;
  ram[34441]  = 1;
  ram[34442]  = 0;
  ram[34443]  = 1;
  ram[34444]  = 1;
  ram[34445]  = 1;
  ram[34446]  = 0;
  ram[34447]  = 1;
  ram[34448]  = 1;
  ram[34449]  = 1;
  ram[34450]  = 1;
  ram[34451]  = 1;
  ram[34452]  = 1;
  ram[34453]  = 0;
  ram[34454]  = 1;
  ram[34455]  = 1;
  ram[34456]  = 1;
  ram[34457]  = 1;
  ram[34458]  = 1;
  ram[34459]  = 1;
  ram[34460]  = 1;
  ram[34461]  = 1;
  ram[34462]  = 0;
  ram[34463]  = 1;
  ram[34464]  = 1;
  ram[34465]  = 1;
  ram[34466]  = 0;
  ram[34467]  = 0;
  ram[34468]  = 1;
  ram[34469]  = 1;
  ram[34470]  = 1;
  ram[34471]  = 1;
  ram[34472]  = 0;
  ram[34473]  = 1;
  ram[34474]  = 1;
  ram[34475]  = 1;
  ram[34476]  = 1;
  ram[34477]  = 1;
  ram[34478]  = 0;
  ram[34479]  = 0;
  ram[34480]  = 1;
  ram[34481]  = 1;
  ram[34482]  = 1;
  ram[34483]  = 1;
  ram[34484]  = 1;
  ram[34485]  = 1;
  ram[34486]  = 1;
  ram[34487]  = 1;
  ram[34488]  = 1;
  ram[34489]  = 1;
  ram[34490]  = 1;
  ram[34491]  = 1;
  ram[34492]  = 1;
  ram[34493]  = 1;
  ram[34494]  = 1;
  ram[34495]  = 1;
  ram[34496]  = 1;
  ram[34497]  = 1;
  ram[34498]  = 1;
  ram[34499]  = 1;
  ram[34500]  = 1;
  ram[34501]  = 1;
  ram[34502]  = 1;
  ram[34503]  = 1;
  ram[34504]  = 1;
  ram[34505]  = 1;
  ram[34506]  = 1;
  ram[34507]  = 1;
  ram[34508]  = 1;
  ram[34509]  = 1;
  ram[34510]  = 1;
  ram[34511]  = 1;
  ram[34512]  = 1;
  ram[34513]  = 1;
  ram[34514]  = 1;
  ram[34515]  = 1;
  ram[34516]  = 0;
  ram[34517]  = 0;
  ram[34518]  = 0;
  ram[34519]  = 1;
  ram[34520]  = 1;
  ram[34521]  = 1;
  ram[34522]  = 1;
  ram[34523]  = 1;
  ram[34524]  = 0;
  ram[34525]  = 1;
  ram[34526]  = 1;
  ram[34527]  = 1;
  ram[34528]  = 1;
  ram[34529]  = 1;
  ram[34530]  = 1;
  ram[34531]  = 0;
  ram[34532]  = 1;
  ram[34533]  = 1;
  ram[34534]  = 0;
  ram[34535]  = 0;
  ram[34536]  = 1;
  ram[34537]  = 1;
  ram[34538]  = 1;
  ram[34539]  = 1;
  ram[34540]  = 1;
  ram[34541]  = 0;
  ram[34542]  = 1;
  ram[34543]  = 1;
  ram[34544]  = 1;
  ram[34545]  = 0;
  ram[34546]  = 1;
  ram[34547]  = 1;
  ram[34548]  = 1;
  ram[34549]  = 1;
  ram[34550]  = 1;
  ram[34551]  = 1;
  ram[34552]  = 1;
  ram[34553]  = 1;
  ram[34554]  = 1;
  ram[34555]  = 1;
  ram[34556]  = 1;
  ram[34557]  = 1;
  ram[34558]  = 0;
  ram[34559]  = 0;
  ram[34560]  = 0;
  ram[34561]  = 1;
  ram[34562]  = 1;
  ram[34563]  = 1;
  ram[34564]  = 1;
  ram[34565]  = 0;
  ram[34566]  = 1;
  ram[34567]  = 1;
  ram[34568]  = 1;
  ram[34569]  = 1;
  ram[34570]  = 1;
  ram[34571]  = 1;
  ram[34572]  = 1;
  ram[34573]  = 1;
  ram[34574]  = 0;
  ram[34575]  = 1;
  ram[34576]  = 1;
  ram[34577]  = 1;
  ram[34578]  = 1;
  ram[34579]  = 1;
  ram[34580]  = 1;
  ram[34581]  = 0;
  ram[34582]  = 1;
  ram[34583]  = 1;
  ram[34584]  = 1;
  ram[34585]  = 0;
  ram[34586]  = 1;
  ram[34587]  = 1;
  ram[34588]  = 1;
  ram[34589]  = 1;
  ram[34590]  = 1;
  ram[34591]  = 0;
  ram[34592]  = 1;
  ram[34593]  = 1;
  ram[34594]  = 1;
  ram[34595]  = 1;
  ram[34596]  = 1;
  ram[34597]  = 0;
  ram[34598]  = 1;
  ram[34599]  = 1;
  ram[34600]  = 1;
  ram[34601]  = 1;
  ram[34602]  = 1;
  ram[34603]  = 1;
  ram[34604]  = 1;
  ram[34605]  = 0;
  ram[34606]  = 0;
  ram[34607]  = 1;
  ram[34608]  = 1;
  ram[34609]  = 0;
  ram[34610]  = 1;
  ram[34611]  = 1;
  ram[34612]  = 1;
  ram[34613]  = 1;
  ram[34614]  = 1;
  ram[34615]  = 1;
  ram[34616]  = 1;
  ram[34617]  = 1;
  ram[34618]  = 1;
  ram[34619]  = 1;
  ram[34620]  = 1;
  ram[34621]  = 1;
  ram[34622]  = 0;
  ram[34623]  = 1;
  ram[34624]  = 1;
  ram[34625]  = 1;
  ram[34626]  = 1;
  ram[34627]  = 1;
  ram[34628]  = 1;
  ram[34629]  = 1;
  ram[34630]  = 0;
  ram[34631]  = 1;
  ram[34632]  = 1;
  ram[34633]  = 1;
  ram[34634]  = 1;
  ram[34635]  = 1;
  ram[34636]  = 0;
  ram[34637]  = 1;
  ram[34638]  = 1;
  ram[34639]  = 1;
  ram[34640]  = 0;
  ram[34641]  = 1;
  ram[34642]  = 1;
  ram[34643]  = 1;
  ram[34644]  = 1;
  ram[34645]  = 1;
  ram[34646]  = 1;
  ram[34647]  = 0;
  ram[34648]  = 1;
  ram[34649]  = 1;
  ram[34650]  = 0;
  ram[34651]  = 1;
  ram[34652]  = 1;
  ram[34653]  = 1;
  ram[34654]  = 0;
  ram[34655]  = 1;
  ram[34656]  = 0;
  ram[34657]  = 1;
  ram[34658]  = 1;
  ram[34659]  = 1;
  ram[34660]  = 0;
  ram[34661]  = 1;
  ram[34662]  = 1;
  ram[34663]  = 1;
  ram[34664]  = 0;
  ram[34665]  = 1;
  ram[34666]  = 1;
  ram[34667]  = 1;
  ram[34668]  = 1;
  ram[34669]  = 1;
  ram[34670]  = 0;
  ram[34671]  = 1;
  ram[34672]  = 1;
  ram[34673]  = 1;
  ram[34674]  = 1;
  ram[34675]  = 1;
  ram[34676]  = 1;
  ram[34677]  = 1;
  ram[34678]  = 1;
  ram[34679]  = 0;
  ram[34680]  = 1;
  ram[34681]  = 1;
  ram[34682]  = 1;
  ram[34683]  = 1;
  ram[34684]  = 1;
  ram[34685]  = 1;
  ram[34686]  = 0;
  ram[34687]  = 1;
  ram[34688]  = 1;
  ram[34689]  = 1;
  ram[34690]  = 0;
  ram[34691]  = 1;
  ram[34692]  = 1;
  ram[34693]  = 1;
  ram[34694]  = 1;
  ram[34695]  = 1;
  ram[34696]  = 0;
  ram[34697]  = 1;
  ram[34698]  = 1;
  ram[34699]  = 1;
  ram[34700]  = 1;
  ram[34701]  = 1;
  ram[34702]  = 1;
  ram[34703]  = 1;
  ram[34704]  = 1;
  ram[34705]  = 0;
  ram[34706]  = 1;
  ram[34707]  = 1;
  ram[34708]  = 1;
  ram[34709]  = 1;
  ram[34710]  = 1;
  ram[34711]  = 0;
  ram[34712]  = 1;
  ram[34713]  = 1;
  ram[34714]  = 1;
  ram[34715]  = 1;
  ram[34716]  = 1;
  ram[34717]  = 0;
  ram[34718]  = 1;
  ram[34719]  = 1;
  ram[34720]  = 0;
  ram[34721]  = 0;
  ram[34722]  = 1;
  ram[34723]  = 1;
  ram[34724]  = 1;
  ram[34725]  = 1;
  ram[34726]  = 1;
  ram[34727]  = 0;
  ram[34728]  = 1;
  ram[34729]  = 1;
  ram[34730]  = 1;
  ram[34731]  = 1;
  ram[34732]  = 1;
  ram[34733]  = 1;
  ram[34734]  = 1;
  ram[34735]  = 0;
  ram[34736]  = 0;
  ram[34737]  = 1;
  ram[34738]  = 1;
  ram[34739]  = 1;
  ram[34740]  = 1;
  ram[34741]  = 1;
  ram[34742]  = 0;
  ram[34743]  = 0;
  ram[34744]  = 1;
  ram[34745]  = 1;
  ram[34746]  = 0;
  ram[34747]  = 1;
  ram[34748]  = 1;
  ram[34749]  = 1;
  ram[34750]  = 1;
  ram[34751]  = 1;
  ram[34752]  = 1;
  ram[34753]  = 0;
  ram[34754]  = 1;
  ram[34755]  = 1;
  ram[34756]  = 1;
  ram[34757]  = 1;
  ram[34758]  = 1;
  ram[34759]  = 1;
  ram[34760]  = 1;
  ram[34761]  = 1;
  ram[34762]  = 0;
  ram[34763]  = 1;
  ram[34764]  = 1;
  ram[34765]  = 1;
  ram[34766]  = 0;
  ram[34767]  = 0;
  ram[34768]  = 1;
  ram[34769]  = 1;
  ram[34770]  = 1;
  ram[34771]  = 1;
  ram[34772]  = 0;
  ram[34773]  = 1;
  ram[34774]  = 1;
  ram[34775]  = 1;
  ram[34776]  = 1;
  ram[34777]  = 1;
  ram[34778]  = 1;
  ram[34779]  = 0;
  ram[34780]  = 1;
  ram[34781]  = 1;
  ram[34782]  = 1;
  ram[34783]  = 1;
  ram[34784]  = 1;
  ram[34785]  = 1;
  ram[34786]  = 1;
  ram[34787]  = 1;
  ram[34788]  = 1;
  ram[34789]  = 1;
  ram[34790]  = 1;
  ram[34791]  = 1;
  ram[34792]  = 1;
  ram[34793]  = 1;
  ram[34794]  = 1;
  ram[34795]  = 1;
  ram[34796]  = 1;
  ram[34797]  = 1;
  ram[34798]  = 1;
  ram[34799]  = 1;
  ram[34800]  = 1;
  ram[34801]  = 1;
  ram[34802]  = 1;
  ram[34803]  = 1;
  ram[34804]  = 1;
  ram[34805]  = 1;
  ram[34806]  = 1;
  ram[34807]  = 1;
  ram[34808]  = 1;
  ram[34809]  = 1;
  ram[34810]  = 1;
  ram[34811]  = 1;
  ram[34812]  = 1;
  ram[34813]  = 1;
  ram[34814]  = 1;
  ram[34815]  = 1;
  ram[34816]  = 0;
  ram[34817]  = 0;
  ram[34818]  = 1;
  ram[34819]  = 1;
  ram[34820]  = 1;
  ram[34821]  = 1;
  ram[34822]  = 1;
  ram[34823]  = 0;
  ram[34824]  = 0;
  ram[34825]  = 1;
  ram[34826]  = 1;
  ram[34827]  = 1;
  ram[34828]  = 1;
  ram[34829]  = 1;
  ram[34830]  = 1;
  ram[34831]  = 0;
  ram[34832]  = 1;
  ram[34833]  = 1;
  ram[34834]  = 0;
  ram[34835]  = 0;
  ram[34836]  = 1;
  ram[34837]  = 1;
  ram[34838]  = 1;
  ram[34839]  = 1;
  ram[34840]  = 1;
  ram[34841]  = 0;
  ram[34842]  = 1;
  ram[34843]  = 1;
  ram[34844]  = 1;
  ram[34845]  = 0;
  ram[34846]  = 1;
  ram[34847]  = 1;
  ram[34848]  = 1;
  ram[34849]  = 1;
  ram[34850]  = 1;
  ram[34851]  = 1;
  ram[34852]  = 1;
  ram[34853]  = 1;
  ram[34854]  = 1;
  ram[34855]  = 1;
  ram[34856]  = 1;
  ram[34857]  = 1;
  ram[34858]  = 1;
  ram[34859]  = 0;
  ram[34860]  = 0;
  ram[34861]  = 0;
  ram[34862]  = 1;
  ram[34863]  = 1;
  ram[34864]  = 1;
  ram[34865]  = 0;
  ram[34866]  = 1;
  ram[34867]  = 1;
  ram[34868]  = 1;
  ram[34869]  = 1;
  ram[34870]  = 1;
  ram[34871]  = 1;
  ram[34872]  = 1;
  ram[34873]  = 1;
  ram[34874]  = 0;
  ram[34875]  = 1;
  ram[34876]  = 1;
  ram[34877]  = 1;
  ram[34878]  = 1;
  ram[34879]  = 1;
  ram[34880]  = 1;
  ram[34881]  = 0;
  ram[34882]  = 1;
  ram[34883]  = 1;
  ram[34884]  = 1;
  ram[34885]  = 0;
  ram[34886]  = 1;
  ram[34887]  = 1;
  ram[34888]  = 1;
  ram[34889]  = 1;
  ram[34890]  = 0;
  ram[34891]  = 0;
  ram[34892]  = 1;
  ram[34893]  = 1;
  ram[34894]  = 1;
  ram[34895]  = 1;
  ram[34896]  = 1;
  ram[34897]  = 0;
  ram[34898]  = 1;
  ram[34899]  = 1;
  ram[34900]  = 1;
  ram[34901]  = 1;
  ram[34902]  = 1;
  ram[34903]  = 1;
  ram[34904]  = 1;
  ram[34905]  = 0;
  ram[34906]  = 0;
  ram[34907]  = 1;
  ram[34908]  = 1;
  ram[34909]  = 0;
  ram[34910]  = 1;
  ram[34911]  = 1;
  ram[34912]  = 1;
  ram[34913]  = 1;
  ram[34914]  = 1;
  ram[34915]  = 1;
  ram[34916]  = 1;
  ram[34917]  = 1;
  ram[34918]  = 1;
  ram[34919]  = 1;
  ram[34920]  = 1;
  ram[34921]  = 1;
  ram[34922]  = 0;
  ram[34923]  = 1;
  ram[34924]  = 1;
  ram[34925]  = 1;
  ram[34926]  = 1;
  ram[34927]  = 1;
  ram[34928]  = 1;
  ram[34929]  = 1;
  ram[34930]  = 0;
  ram[34931]  = 1;
  ram[34932]  = 1;
  ram[34933]  = 1;
  ram[34934]  = 1;
  ram[34935]  = 1;
  ram[34936]  = 0;
  ram[34937]  = 1;
  ram[34938]  = 1;
  ram[34939]  = 1;
  ram[34940]  = 0;
  ram[34941]  = 1;
  ram[34942]  = 1;
  ram[34943]  = 1;
  ram[34944]  = 1;
  ram[34945]  = 1;
  ram[34946]  = 1;
  ram[34947]  = 0;
  ram[34948]  = 1;
  ram[34949]  = 1;
  ram[34950]  = 0;
  ram[34951]  = 1;
  ram[34952]  = 1;
  ram[34953]  = 1;
  ram[34954]  = 0;
  ram[34955]  = 1;
  ram[34956]  = 0;
  ram[34957]  = 1;
  ram[34958]  = 1;
  ram[34959]  = 1;
  ram[34960]  = 0;
  ram[34961]  = 1;
  ram[34962]  = 1;
  ram[34963]  = 1;
  ram[34964]  = 0;
  ram[34965]  = 1;
  ram[34966]  = 1;
  ram[34967]  = 1;
  ram[34968]  = 1;
  ram[34969]  = 1;
  ram[34970]  = 0;
  ram[34971]  = 1;
  ram[34972]  = 1;
  ram[34973]  = 1;
  ram[34974]  = 1;
  ram[34975]  = 1;
  ram[34976]  = 1;
  ram[34977]  = 1;
  ram[34978]  = 0;
  ram[34979]  = 0;
  ram[34980]  = 1;
  ram[34981]  = 1;
  ram[34982]  = 1;
  ram[34983]  = 1;
  ram[34984]  = 1;
  ram[34985]  = 1;
  ram[34986]  = 0;
  ram[34987]  = 1;
  ram[34988]  = 1;
  ram[34989]  = 1;
  ram[34990]  = 0;
  ram[34991]  = 1;
  ram[34992]  = 1;
  ram[34993]  = 1;
  ram[34994]  = 1;
  ram[34995]  = 1;
  ram[34996]  = 0;
  ram[34997]  = 1;
  ram[34998]  = 1;
  ram[34999]  = 1;
  ram[35000]  = 1;
  ram[35001]  = 1;
  ram[35002]  = 1;
  ram[35003]  = 1;
  ram[35004]  = 1;
  ram[35005]  = 0;
  ram[35006]  = 1;
  ram[35007]  = 1;
  ram[35008]  = 1;
  ram[35009]  = 1;
  ram[35010]  = 1;
  ram[35011]  = 0;
  ram[35012]  = 1;
  ram[35013]  = 1;
  ram[35014]  = 1;
  ram[35015]  = 1;
  ram[35016]  = 1;
  ram[35017]  = 0;
  ram[35018]  = 1;
  ram[35019]  = 1;
  ram[35020]  = 0;
  ram[35021]  = 0;
  ram[35022]  = 1;
  ram[35023]  = 1;
  ram[35024]  = 1;
  ram[35025]  = 1;
  ram[35026]  = 1;
  ram[35027]  = 0;
  ram[35028]  = 1;
  ram[35029]  = 1;
  ram[35030]  = 1;
  ram[35031]  = 1;
  ram[35032]  = 1;
  ram[35033]  = 1;
  ram[35034]  = 1;
  ram[35035]  = 0;
  ram[35036]  = 0;
  ram[35037]  = 1;
  ram[35038]  = 1;
  ram[35039]  = 1;
  ram[35040]  = 1;
  ram[35041]  = 1;
  ram[35042]  = 0;
  ram[35043]  = 0;
  ram[35044]  = 1;
  ram[35045]  = 1;
  ram[35046]  = 0;
  ram[35047]  = 1;
  ram[35048]  = 1;
  ram[35049]  = 1;
  ram[35050]  = 1;
  ram[35051]  = 1;
  ram[35052]  = 1;
  ram[35053]  = 0;
  ram[35054]  = 1;
  ram[35055]  = 1;
  ram[35056]  = 1;
  ram[35057]  = 1;
  ram[35058]  = 1;
  ram[35059]  = 1;
  ram[35060]  = 1;
  ram[35061]  = 1;
  ram[35062]  = 0;
  ram[35063]  = 1;
  ram[35064]  = 1;
  ram[35065]  = 1;
  ram[35066]  = 0;
  ram[35067]  = 1;
  ram[35068]  = 1;
  ram[35069]  = 1;
  ram[35070]  = 1;
  ram[35071]  = 1;
  ram[35072]  = 0;
  ram[35073]  = 1;
  ram[35074]  = 1;
  ram[35075]  = 1;
  ram[35076]  = 1;
  ram[35077]  = 1;
  ram[35078]  = 1;
  ram[35079]  = 0;
  ram[35080]  = 1;
  ram[35081]  = 1;
  ram[35082]  = 1;
  ram[35083]  = 1;
  ram[35084]  = 1;
  ram[35085]  = 1;
  ram[35086]  = 1;
  ram[35087]  = 1;
  ram[35088]  = 1;
  ram[35089]  = 1;
  ram[35090]  = 1;
  ram[35091]  = 1;
  ram[35092]  = 1;
  ram[35093]  = 1;
  ram[35094]  = 1;
  ram[35095]  = 1;
  ram[35096]  = 1;
  ram[35097]  = 1;
  ram[35098]  = 1;
  ram[35099]  = 1;
  ram[35100]  = 1;
  ram[35101]  = 1;
  ram[35102]  = 1;
  ram[35103]  = 1;
  ram[35104]  = 1;
  ram[35105]  = 1;
  ram[35106]  = 1;
  ram[35107]  = 1;
  ram[35108]  = 1;
  ram[35109]  = 1;
  ram[35110]  = 1;
  ram[35111]  = 1;
  ram[35112]  = 1;
  ram[35113]  = 1;
  ram[35114]  = 1;
  ram[35115]  = 1;
  ram[35116]  = 1;
  ram[35117]  = 0;
  ram[35118]  = 1;
  ram[35119]  = 1;
  ram[35120]  = 1;
  ram[35121]  = 1;
  ram[35122]  = 1;
  ram[35123]  = 0;
  ram[35124]  = 0;
  ram[35125]  = 1;
  ram[35126]  = 1;
  ram[35127]  = 1;
  ram[35128]  = 1;
  ram[35129]  = 1;
  ram[35130]  = 1;
  ram[35131]  = 0;
  ram[35132]  = 1;
  ram[35133]  = 1;
  ram[35134]  = 0;
  ram[35135]  = 0;
  ram[35136]  = 1;
  ram[35137]  = 1;
  ram[35138]  = 1;
  ram[35139]  = 1;
  ram[35140]  = 1;
  ram[35141]  = 0;
  ram[35142]  = 1;
  ram[35143]  = 1;
  ram[35144]  = 1;
  ram[35145]  = 0;
  ram[35146]  = 1;
  ram[35147]  = 1;
  ram[35148]  = 1;
  ram[35149]  = 1;
  ram[35150]  = 1;
  ram[35151]  = 1;
  ram[35152]  = 1;
  ram[35153]  = 1;
  ram[35154]  = 1;
  ram[35155]  = 1;
  ram[35156]  = 1;
  ram[35157]  = 1;
  ram[35158]  = 1;
  ram[35159]  = 1;
  ram[35160]  = 1;
  ram[35161]  = 0;
  ram[35162]  = 0;
  ram[35163]  = 1;
  ram[35164]  = 1;
  ram[35165]  = 0;
  ram[35166]  = 1;
  ram[35167]  = 1;
  ram[35168]  = 1;
  ram[35169]  = 1;
  ram[35170]  = 1;
  ram[35171]  = 1;
  ram[35172]  = 1;
  ram[35173]  = 0;
  ram[35174]  = 0;
  ram[35175]  = 1;
  ram[35176]  = 1;
  ram[35177]  = 1;
  ram[35178]  = 1;
  ram[35179]  = 1;
  ram[35180]  = 1;
  ram[35181]  = 0;
  ram[35182]  = 1;
  ram[35183]  = 1;
  ram[35184]  = 1;
  ram[35185]  = 0;
  ram[35186]  = 1;
  ram[35187]  = 1;
  ram[35188]  = 1;
  ram[35189]  = 1;
  ram[35190]  = 0;
  ram[35191]  = 0;
  ram[35192]  = 1;
  ram[35193]  = 1;
  ram[35194]  = 1;
  ram[35195]  = 1;
  ram[35196]  = 1;
  ram[35197]  = 0;
  ram[35198]  = 1;
  ram[35199]  = 1;
  ram[35200]  = 1;
  ram[35201]  = 1;
  ram[35202]  = 1;
  ram[35203]  = 1;
  ram[35204]  = 1;
  ram[35205]  = 0;
  ram[35206]  = 0;
  ram[35207]  = 1;
  ram[35208]  = 1;
  ram[35209]  = 0;
  ram[35210]  = 0;
  ram[35211]  = 0;
  ram[35212]  = 1;
  ram[35213]  = 1;
  ram[35214]  = 1;
  ram[35215]  = 1;
  ram[35216]  = 1;
  ram[35217]  = 1;
  ram[35218]  = 1;
  ram[35219]  = 1;
  ram[35220]  = 1;
  ram[35221]  = 1;
  ram[35222]  = 0;
  ram[35223]  = 0;
  ram[35224]  = 1;
  ram[35225]  = 1;
  ram[35226]  = 1;
  ram[35227]  = 1;
  ram[35228]  = 1;
  ram[35229]  = 1;
  ram[35230]  = 0;
  ram[35231]  = 1;
  ram[35232]  = 1;
  ram[35233]  = 1;
  ram[35234]  = 1;
  ram[35235]  = 1;
  ram[35236]  = 0;
  ram[35237]  = 1;
  ram[35238]  = 1;
  ram[35239]  = 0;
  ram[35240]  = 0;
  ram[35241]  = 1;
  ram[35242]  = 1;
  ram[35243]  = 1;
  ram[35244]  = 1;
  ram[35245]  = 1;
  ram[35246]  = 1;
  ram[35247]  = 0;
  ram[35248]  = 1;
  ram[35249]  = 1;
  ram[35250]  = 0;
  ram[35251]  = 0;
  ram[35252]  = 1;
  ram[35253]  = 1;
  ram[35254]  = 0;
  ram[35255]  = 1;
  ram[35256]  = 0;
  ram[35257]  = 1;
  ram[35258]  = 1;
  ram[35259]  = 1;
  ram[35260]  = 0;
  ram[35261]  = 1;
  ram[35262]  = 1;
  ram[35263]  = 1;
  ram[35264]  = 0;
  ram[35265]  = 1;
  ram[35266]  = 1;
  ram[35267]  = 1;
  ram[35268]  = 1;
  ram[35269]  = 1;
  ram[35270]  = 0;
  ram[35271]  = 1;
  ram[35272]  = 1;
  ram[35273]  = 1;
  ram[35274]  = 1;
  ram[35275]  = 1;
  ram[35276]  = 1;
  ram[35277]  = 1;
  ram[35278]  = 0;
  ram[35279]  = 0;
  ram[35280]  = 1;
  ram[35281]  = 1;
  ram[35282]  = 1;
  ram[35283]  = 1;
  ram[35284]  = 1;
  ram[35285]  = 1;
  ram[35286]  = 0;
  ram[35287]  = 1;
  ram[35288]  = 1;
  ram[35289]  = 1;
  ram[35290]  = 0;
  ram[35291]  = 1;
  ram[35292]  = 1;
  ram[35293]  = 1;
  ram[35294]  = 1;
  ram[35295]  = 1;
  ram[35296]  = 0;
  ram[35297]  = 1;
  ram[35298]  = 1;
  ram[35299]  = 1;
  ram[35300]  = 1;
  ram[35301]  = 1;
  ram[35302]  = 1;
  ram[35303]  = 1;
  ram[35304]  = 1;
  ram[35305]  = 0;
  ram[35306]  = 1;
  ram[35307]  = 1;
  ram[35308]  = 1;
  ram[35309]  = 1;
  ram[35310]  = 1;
  ram[35311]  = 0;
  ram[35312]  = 1;
  ram[35313]  = 1;
  ram[35314]  = 1;
  ram[35315]  = 1;
  ram[35316]  = 1;
  ram[35317]  = 0;
  ram[35318]  = 1;
  ram[35319]  = 1;
  ram[35320]  = 0;
  ram[35321]  = 0;
  ram[35322]  = 1;
  ram[35323]  = 1;
  ram[35324]  = 1;
  ram[35325]  = 1;
  ram[35326]  = 1;
  ram[35327]  = 0;
  ram[35328]  = 1;
  ram[35329]  = 1;
  ram[35330]  = 1;
  ram[35331]  = 1;
  ram[35332]  = 1;
  ram[35333]  = 1;
  ram[35334]  = 1;
  ram[35335]  = 0;
  ram[35336]  = 0;
  ram[35337]  = 1;
  ram[35338]  = 1;
  ram[35339]  = 1;
  ram[35340]  = 1;
  ram[35341]  = 1;
  ram[35342]  = 0;
  ram[35343]  = 0;
  ram[35344]  = 1;
  ram[35345]  = 1;
  ram[35346]  = 0;
  ram[35347]  = 1;
  ram[35348]  = 1;
  ram[35349]  = 1;
  ram[35350]  = 1;
  ram[35351]  = 1;
  ram[35352]  = 1;
  ram[35353]  = 0;
  ram[35354]  = 1;
  ram[35355]  = 1;
  ram[35356]  = 1;
  ram[35357]  = 1;
  ram[35358]  = 1;
  ram[35359]  = 0;
  ram[35360]  = 0;
  ram[35361]  = 0;
  ram[35362]  = 0;
  ram[35363]  = 1;
  ram[35364]  = 1;
  ram[35365]  = 1;
  ram[35366]  = 0;
  ram[35367]  = 1;
  ram[35368]  = 1;
  ram[35369]  = 1;
  ram[35370]  = 1;
  ram[35371]  = 1;
  ram[35372]  = 0;
  ram[35373]  = 1;
  ram[35374]  = 1;
  ram[35375]  = 1;
  ram[35376]  = 1;
  ram[35377]  = 1;
  ram[35378]  = 1;
  ram[35379]  = 0;
  ram[35380]  = 1;
  ram[35381]  = 1;
  ram[35382]  = 1;
  ram[35383]  = 1;
  ram[35384]  = 1;
  ram[35385]  = 1;
  ram[35386]  = 1;
  ram[35387]  = 1;
  ram[35388]  = 1;
  ram[35389]  = 1;
  ram[35390]  = 1;
  ram[35391]  = 1;
  ram[35392]  = 1;
  ram[35393]  = 1;
  ram[35394]  = 1;
  ram[35395]  = 1;
  ram[35396]  = 1;
  ram[35397]  = 1;
  ram[35398]  = 1;
  ram[35399]  = 1;
  ram[35400]  = 1;
  ram[35401]  = 1;
  ram[35402]  = 1;
  ram[35403]  = 1;
  ram[35404]  = 1;
  ram[35405]  = 1;
  ram[35406]  = 1;
  ram[35407]  = 1;
  ram[35408]  = 1;
  ram[35409]  = 1;
  ram[35410]  = 1;
  ram[35411]  = 1;
  ram[35412]  = 1;
  ram[35413]  = 1;
  ram[35414]  = 1;
  ram[35415]  = 1;
  ram[35416]  = 1;
  ram[35417]  = 0;
  ram[35418]  = 1;
  ram[35419]  = 1;
  ram[35420]  = 1;
  ram[35421]  = 1;
  ram[35422]  = 1;
  ram[35423]  = 0;
  ram[35424]  = 0;
  ram[35425]  = 1;
  ram[35426]  = 1;
  ram[35427]  = 1;
  ram[35428]  = 1;
  ram[35429]  = 1;
  ram[35430]  = 1;
  ram[35431]  = 0;
  ram[35432]  = 1;
  ram[35433]  = 1;
  ram[35434]  = 0;
  ram[35435]  = 0;
  ram[35436]  = 1;
  ram[35437]  = 1;
  ram[35438]  = 1;
  ram[35439]  = 1;
  ram[35440]  = 1;
  ram[35441]  = 0;
  ram[35442]  = 1;
  ram[35443]  = 1;
  ram[35444]  = 1;
  ram[35445]  = 0;
  ram[35446]  = 1;
  ram[35447]  = 1;
  ram[35448]  = 1;
  ram[35449]  = 1;
  ram[35450]  = 1;
  ram[35451]  = 1;
  ram[35452]  = 1;
  ram[35453]  = 1;
  ram[35454]  = 1;
  ram[35455]  = 1;
  ram[35456]  = 1;
  ram[35457]  = 1;
  ram[35458]  = 1;
  ram[35459]  = 1;
  ram[35460]  = 1;
  ram[35461]  = 1;
  ram[35462]  = 0;
  ram[35463]  = 1;
  ram[35464]  = 1;
  ram[35465]  = 0;
  ram[35466]  = 1;
  ram[35467]  = 1;
  ram[35468]  = 1;
  ram[35469]  = 1;
  ram[35470]  = 1;
  ram[35471]  = 1;
  ram[35472]  = 1;
  ram[35473]  = 0;
  ram[35474]  = 0;
  ram[35475]  = 1;
  ram[35476]  = 1;
  ram[35477]  = 1;
  ram[35478]  = 1;
  ram[35479]  = 1;
  ram[35480]  = 1;
  ram[35481]  = 0;
  ram[35482]  = 1;
  ram[35483]  = 1;
  ram[35484]  = 1;
  ram[35485]  = 0;
  ram[35486]  = 1;
  ram[35487]  = 1;
  ram[35488]  = 1;
  ram[35489]  = 1;
  ram[35490]  = 0;
  ram[35491]  = 0;
  ram[35492]  = 0;
  ram[35493]  = 0;
  ram[35494]  = 0;
  ram[35495]  = 0;
  ram[35496]  = 0;
  ram[35497]  = 0;
  ram[35498]  = 1;
  ram[35499]  = 1;
  ram[35500]  = 1;
  ram[35501]  = 1;
  ram[35502]  = 1;
  ram[35503]  = 1;
  ram[35504]  = 1;
  ram[35505]  = 0;
  ram[35506]  = 0;
  ram[35507]  = 1;
  ram[35508]  = 1;
  ram[35509]  = 1;
  ram[35510]  = 0;
  ram[35511]  = 0;
  ram[35512]  = 0;
  ram[35513]  = 1;
  ram[35514]  = 1;
  ram[35515]  = 1;
  ram[35516]  = 1;
  ram[35517]  = 1;
  ram[35518]  = 1;
  ram[35519]  = 1;
  ram[35520]  = 1;
  ram[35521]  = 1;
  ram[35522]  = 1;
  ram[35523]  = 0;
  ram[35524]  = 0;
  ram[35525]  = 0;
  ram[35526]  = 1;
  ram[35527]  = 1;
  ram[35528]  = 1;
  ram[35529]  = 1;
  ram[35530]  = 0;
  ram[35531]  = 1;
  ram[35532]  = 1;
  ram[35533]  = 1;
  ram[35534]  = 1;
  ram[35535]  = 1;
  ram[35536]  = 0;
  ram[35537]  = 1;
  ram[35538]  = 1;
  ram[35539]  = 0;
  ram[35540]  = 0;
  ram[35541]  = 1;
  ram[35542]  = 1;
  ram[35543]  = 1;
  ram[35544]  = 1;
  ram[35545]  = 1;
  ram[35546]  = 1;
  ram[35547]  = 0;
  ram[35548]  = 1;
  ram[35549]  = 1;
  ram[35550]  = 1;
  ram[35551]  = 0;
  ram[35552]  = 1;
  ram[35553]  = 1;
  ram[35554]  = 0;
  ram[35555]  = 1;
  ram[35556]  = 0;
  ram[35557]  = 1;
  ram[35558]  = 1;
  ram[35559]  = 0;
  ram[35560]  = 0;
  ram[35561]  = 1;
  ram[35562]  = 1;
  ram[35563]  = 1;
  ram[35564]  = 0;
  ram[35565]  = 1;
  ram[35566]  = 1;
  ram[35567]  = 1;
  ram[35568]  = 1;
  ram[35569]  = 1;
  ram[35570]  = 0;
  ram[35571]  = 1;
  ram[35572]  = 1;
  ram[35573]  = 1;
  ram[35574]  = 1;
  ram[35575]  = 1;
  ram[35576]  = 1;
  ram[35577]  = 1;
  ram[35578]  = 0;
  ram[35579]  = 0;
  ram[35580]  = 1;
  ram[35581]  = 1;
  ram[35582]  = 1;
  ram[35583]  = 1;
  ram[35584]  = 1;
  ram[35585]  = 1;
  ram[35586]  = 0;
  ram[35587]  = 1;
  ram[35588]  = 1;
  ram[35589]  = 1;
  ram[35590]  = 0;
  ram[35591]  = 1;
  ram[35592]  = 1;
  ram[35593]  = 1;
  ram[35594]  = 1;
  ram[35595]  = 1;
  ram[35596]  = 0;
  ram[35597]  = 1;
  ram[35598]  = 1;
  ram[35599]  = 1;
  ram[35600]  = 1;
  ram[35601]  = 1;
  ram[35602]  = 1;
  ram[35603]  = 1;
  ram[35604]  = 1;
  ram[35605]  = 0;
  ram[35606]  = 1;
  ram[35607]  = 1;
  ram[35608]  = 1;
  ram[35609]  = 1;
  ram[35610]  = 1;
  ram[35611]  = 0;
  ram[35612]  = 1;
  ram[35613]  = 1;
  ram[35614]  = 1;
  ram[35615]  = 1;
  ram[35616]  = 1;
  ram[35617]  = 0;
  ram[35618]  = 1;
  ram[35619]  = 1;
  ram[35620]  = 0;
  ram[35621]  = 0;
  ram[35622]  = 0;
  ram[35623]  = 0;
  ram[35624]  = 0;
  ram[35625]  = 0;
  ram[35626]  = 0;
  ram[35627]  = 0;
  ram[35628]  = 1;
  ram[35629]  = 1;
  ram[35630]  = 1;
  ram[35631]  = 1;
  ram[35632]  = 1;
  ram[35633]  = 1;
  ram[35634]  = 1;
  ram[35635]  = 0;
  ram[35636]  = 0;
  ram[35637]  = 1;
  ram[35638]  = 1;
  ram[35639]  = 1;
  ram[35640]  = 1;
  ram[35641]  = 1;
  ram[35642]  = 1;
  ram[35643]  = 0;
  ram[35644]  = 1;
  ram[35645]  = 1;
  ram[35646]  = 0;
  ram[35647]  = 1;
  ram[35648]  = 1;
  ram[35649]  = 1;
  ram[35650]  = 1;
  ram[35651]  = 1;
  ram[35652]  = 1;
  ram[35653]  = 0;
  ram[35654]  = 1;
  ram[35655]  = 1;
  ram[35656]  = 1;
  ram[35657]  = 0;
  ram[35658]  = 0;
  ram[35659]  = 0;
  ram[35660]  = 0;
  ram[35661]  = 0;
  ram[35662]  = 0;
  ram[35663]  = 1;
  ram[35664]  = 1;
  ram[35665]  = 1;
  ram[35666]  = 0;
  ram[35667]  = 1;
  ram[35668]  = 1;
  ram[35669]  = 1;
  ram[35670]  = 1;
  ram[35671]  = 1;
  ram[35672]  = 0;
  ram[35673]  = 1;
  ram[35674]  = 1;
  ram[35675]  = 1;
  ram[35676]  = 1;
  ram[35677]  = 1;
  ram[35678]  = 1;
  ram[35679]  = 0;
  ram[35680]  = 1;
  ram[35681]  = 1;
  ram[35682]  = 1;
  ram[35683]  = 1;
  ram[35684]  = 1;
  ram[35685]  = 1;
  ram[35686]  = 1;
  ram[35687]  = 1;
  ram[35688]  = 1;
  ram[35689]  = 1;
  ram[35690]  = 1;
  ram[35691]  = 1;
  ram[35692]  = 1;
  ram[35693]  = 1;
  ram[35694]  = 1;
  ram[35695]  = 1;
  ram[35696]  = 1;
  ram[35697]  = 1;
  ram[35698]  = 1;
  ram[35699]  = 1;
  ram[35700]  = 1;
  ram[35701]  = 1;
  ram[35702]  = 1;
  ram[35703]  = 1;
  ram[35704]  = 1;
  ram[35705]  = 1;
  ram[35706]  = 1;
  ram[35707]  = 1;
  ram[35708]  = 1;
  ram[35709]  = 1;
  ram[35710]  = 1;
  ram[35711]  = 1;
  ram[35712]  = 1;
  ram[35713]  = 1;
  ram[35714]  = 1;
  ram[35715]  = 1;
  ram[35716]  = 1;
  ram[35717]  = 0;
  ram[35718]  = 1;
  ram[35719]  = 1;
  ram[35720]  = 1;
  ram[35721]  = 1;
  ram[35722]  = 1;
  ram[35723]  = 0;
  ram[35724]  = 0;
  ram[35725]  = 1;
  ram[35726]  = 1;
  ram[35727]  = 1;
  ram[35728]  = 1;
  ram[35729]  = 1;
  ram[35730]  = 1;
  ram[35731]  = 0;
  ram[35732]  = 1;
  ram[35733]  = 1;
  ram[35734]  = 0;
  ram[35735]  = 0;
  ram[35736]  = 1;
  ram[35737]  = 1;
  ram[35738]  = 1;
  ram[35739]  = 1;
  ram[35740]  = 1;
  ram[35741]  = 0;
  ram[35742]  = 1;
  ram[35743]  = 1;
  ram[35744]  = 1;
  ram[35745]  = 0;
  ram[35746]  = 1;
  ram[35747]  = 1;
  ram[35748]  = 1;
  ram[35749]  = 1;
  ram[35750]  = 1;
  ram[35751]  = 1;
  ram[35752]  = 1;
  ram[35753]  = 1;
  ram[35754]  = 1;
  ram[35755]  = 1;
  ram[35756]  = 1;
  ram[35757]  = 1;
  ram[35758]  = 1;
  ram[35759]  = 1;
  ram[35760]  = 1;
  ram[35761]  = 1;
  ram[35762]  = 0;
  ram[35763]  = 1;
  ram[35764]  = 1;
  ram[35765]  = 0;
  ram[35766]  = 1;
  ram[35767]  = 1;
  ram[35768]  = 1;
  ram[35769]  = 1;
  ram[35770]  = 1;
  ram[35771]  = 1;
  ram[35772]  = 1;
  ram[35773]  = 0;
  ram[35774]  = 0;
  ram[35775]  = 1;
  ram[35776]  = 1;
  ram[35777]  = 1;
  ram[35778]  = 1;
  ram[35779]  = 1;
  ram[35780]  = 1;
  ram[35781]  = 0;
  ram[35782]  = 1;
  ram[35783]  = 1;
  ram[35784]  = 1;
  ram[35785]  = 0;
  ram[35786]  = 1;
  ram[35787]  = 1;
  ram[35788]  = 1;
  ram[35789]  = 1;
  ram[35790]  = 0;
  ram[35791]  = 0;
  ram[35792]  = 1;
  ram[35793]  = 1;
  ram[35794]  = 1;
  ram[35795]  = 1;
  ram[35796]  = 1;
  ram[35797]  = 1;
  ram[35798]  = 1;
  ram[35799]  = 1;
  ram[35800]  = 1;
  ram[35801]  = 1;
  ram[35802]  = 1;
  ram[35803]  = 1;
  ram[35804]  = 1;
  ram[35805]  = 0;
  ram[35806]  = 0;
  ram[35807]  = 1;
  ram[35808]  = 1;
  ram[35809]  = 1;
  ram[35810]  = 1;
  ram[35811]  = 1;
  ram[35812]  = 0;
  ram[35813]  = 0;
  ram[35814]  = 1;
  ram[35815]  = 1;
  ram[35816]  = 1;
  ram[35817]  = 1;
  ram[35818]  = 1;
  ram[35819]  = 1;
  ram[35820]  = 1;
  ram[35821]  = 1;
  ram[35822]  = 1;
  ram[35823]  = 1;
  ram[35824]  = 0;
  ram[35825]  = 0;
  ram[35826]  = 0;
  ram[35827]  = 1;
  ram[35828]  = 1;
  ram[35829]  = 1;
  ram[35830]  = 0;
  ram[35831]  = 1;
  ram[35832]  = 1;
  ram[35833]  = 1;
  ram[35834]  = 1;
  ram[35835]  = 1;
  ram[35836]  = 0;
  ram[35837]  = 1;
  ram[35838]  = 1;
  ram[35839]  = 0;
  ram[35840]  = 0;
  ram[35841]  = 1;
  ram[35842]  = 1;
  ram[35843]  = 1;
  ram[35844]  = 1;
  ram[35845]  = 1;
  ram[35846]  = 1;
  ram[35847]  = 0;
  ram[35848]  = 1;
  ram[35849]  = 1;
  ram[35850]  = 1;
  ram[35851]  = 0;
  ram[35852]  = 1;
  ram[35853]  = 0;
  ram[35854]  = 0;
  ram[35855]  = 1;
  ram[35856]  = 1;
  ram[35857]  = 0;
  ram[35858]  = 1;
  ram[35859]  = 0;
  ram[35860]  = 1;
  ram[35861]  = 1;
  ram[35862]  = 1;
  ram[35863]  = 1;
  ram[35864]  = 0;
  ram[35865]  = 1;
  ram[35866]  = 1;
  ram[35867]  = 1;
  ram[35868]  = 1;
  ram[35869]  = 1;
  ram[35870]  = 0;
  ram[35871]  = 1;
  ram[35872]  = 1;
  ram[35873]  = 1;
  ram[35874]  = 1;
  ram[35875]  = 1;
  ram[35876]  = 1;
  ram[35877]  = 1;
  ram[35878]  = 0;
  ram[35879]  = 0;
  ram[35880]  = 1;
  ram[35881]  = 1;
  ram[35882]  = 1;
  ram[35883]  = 1;
  ram[35884]  = 1;
  ram[35885]  = 1;
  ram[35886]  = 0;
  ram[35887]  = 1;
  ram[35888]  = 1;
  ram[35889]  = 1;
  ram[35890]  = 0;
  ram[35891]  = 1;
  ram[35892]  = 1;
  ram[35893]  = 1;
  ram[35894]  = 1;
  ram[35895]  = 1;
  ram[35896]  = 0;
  ram[35897]  = 1;
  ram[35898]  = 1;
  ram[35899]  = 1;
  ram[35900]  = 1;
  ram[35901]  = 1;
  ram[35902]  = 1;
  ram[35903]  = 1;
  ram[35904]  = 1;
  ram[35905]  = 0;
  ram[35906]  = 1;
  ram[35907]  = 1;
  ram[35908]  = 1;
  ram[35909]  = 1;
  ram[35910]  = 1;
  ram[35911]  = 0;
  ram[35912]  = 1;
  ram[35913]  = 1;
  ram[35914]  = 1;
  ram[35915]  = 1;
  ram[35916]  = 1;
  ram[35917]  = 0;
  ram[35918]  = 1;
  ram[35919]  = 1;
  ram[35920]  = 0;
  ram[35921]  = 0;
  ram[35922]  = 1;
  ram[35923]  = 1;
  ram[35924]  = 1;
  ram[35925]  = 1;
  ram[35926]  = 1;
  ram[35927]  = 1;
  ram[35928]  = 1;
  ram[35929]  = 1;
  ram[35930]  = 1;
  ram[35931]  = 1;
  ram[35932]  = 1;
  ram[35933]  = 1;
  ram[35934]  = 1;
  ram[35935]  = 0;
  ram[35936]  = 0;
  ram[35937]  = 1;
  ram[35938]  = 1;
  ram[35939]  = 1;
  ram[35940]  = 1;
  ram[35941]  = 1;
  ram[35942]  = 0;
  ram[35943]  = 0;
  ram[35944]  = 1;
  ram[35945]  = 1;
  ram[35946]  = 0;
  ram[35947]  = 1;
  ram[35948]  = 1;
  ram[35949]  = 1;
  ram[35950]  = 1;
  ram[35951]  = 1;
  ram[35952]  = 1;
  ram[35953]  = 0;
  ram[35954]  = 1;
  ram[35955]  = 1;
  ram[35956]  = 1;
  ram[35957]  = 0;
  ram[35958]  = 1;
  ram[35959]  = 1;
  ram[35960]  = 1;
  ram[35961]  = 1;
  ram[35962]  = 0;
  ram[35963]  = 1;
  ram[35964]  = 1;
  ram[35965]  = 1;
  ram[35966]  = 0;
  ram[35967]  = 1;
  ram[35968]  = 1;
  ram[35969]  = 1;
  ram[35970]  = 1;
  ram[35971]  = 1;
  ram[35972]  = 0;
  ram[35973]  = 1;
  ram[35974]  = 1;
  ram[35975]  = 1;
  ram[35976]  = 1;
  ram[35977]  = 1;
  ram[35978]  = 1;
  ram[35979]  = 0;
  ram[35980]  = 1;
  ram[35981]  = 1;
  ram[35982]  = 1;
  ram[35983]  = 1;
  ram[35984]  = 1;
  ram[35985]  = 1;
  ram[35986]  = 1;
  ram[35987]  = 1;
  ram[35988]  = 1;
  ram[35989]  = 1;
  ram[35990]  = 1;
  ram[35991]  = 1;
  ram[35992]  = 1;
  ram[35993]  = 1;
  ram[35994]  = 1;
  ram[35995]  = 1;
  ram[35996]  = 1;
  ram[35997]  = 1;
  ram[35998]  = 1;
  ram[35999]  = 1;
  ram[36000]  = 1;
  ram[36001]  = 1;
  ram[36002]  = 1;
  ram[36003]  = 1;
  ram[36004]  = 1;
  ram[36005]  = 1;
  ram[36006]  = 1;
  ram[36007]  = 1;
  ram[36008]  = 1;
  ram[36009]  = 1;
  ram[36010]  = 1;
  ram[36011]  = 1;
  ram[36012]  = 1;
  ram[36013]  = 1;
  ram[36014]  = 1;
  ram[36015]  = 1;
  ram[36016]  = 1;
  ram[36017]  = 0;
  ram[36018]  = 1;
  ram[36019]  = 1;
  ram[36020]  = 1;
  ram[36021]  = 1;
  ram[36022]  = 1;
  ram[36023]  = 0;
  ram[36024]  = 0;
  ram[36025]  = 1;
  ram[36026]  = 1;
  ram[36027]  = 1;
  ram[36028]  = 1;
  ram[36029]  = 1;
  ram[36030]  = 1;
  ram[36031]  = 0;
  ram[36032]  = 1;
  ram[36033]  = 1;
  ram[36034]  = 0;
  ram[36035]  = 0;
  ram[36036]  = 1;
  ram[36037]  = 1;
  ram[36038]  = 1;
  ram[36039]  = 1;
  ram[36040]  = 1;
  ram[36041]  = 0;
  ram[36042]  = 1;
  ram[36043]  = 1;
  ram[36044]  = 1;
  ram[36045]  = 0;
  ram[36046]  = 1;
  ram[36047]  = 1;
  ram[36048]  = 1;
  ram[36049]  = 1;
  ram[36050]  = 1;
  ram[36051]  = 1;
  ram[36052]  = 1;
  ram[36053]  = 1;
  ram[36054]  = 1;
  ram[36055]  = 1;
  ram[36056]  = 1;
  ram[36057]  = 1;
  ram[36058]  = 1;
  ram[36059]  = 1;
  ram[36060]  = 1;
  ram[36061]  = 1;
  ram[36062]  = 0;
  ram[36063]  = 1;
  ram[36064]  = 1;
  ram[36065]  = 0;
  ram[36066]  = 1;
  ram[36067]  = 1;
  ram[36068]  = 1;
  ram[36069]  = 1;
  ram[36070]  = 1;
  ram[36071]  = 1;
  ram[36072]  = 1;
  ram[36073]  = 0;
  ram[36074]  = 0;
  ram[36075]  = 1;
  ram[36076]  = 1;
  ram[36077]  = 1;
  ram[36078]  = 1;
  ram[36079]  = 1;
  ram[36080]  = 1;
  ram[36081]  = 0;
  ram[36082]  = 1;
  ram[36083]  = 1;
  ram[36084]  = 1;
  ram[36085]  = 0;
  ram[36086]  = 1;
  ram[36087]  = 1;
  ram[36088]  = 1;
  ram[36089]  = 1;
  ram[36090]  = 0;
  ram[36091]  = 0;
  ram[36092]  = 1;
  ram[36093]  = 1;
  ram[36094]  = 1;
  ram[36095]  = 1;
  ram[36096]  = 1;
  ram[36097]  = 1;
  ram[36098]  = 1;
  ram[36099]  = 1;
  ram[36100]  = 1;
  ram[36101]  = 1;
  ram[36102]  = 1;
  ram[36103]  = 1;
  ram[36104]  = 1;
  ram[36105]  = 0;
  ram[36106]  = 0;
  ram[36107]  = 1;
  ram[36108]  = 1;
  ram[36109]  = 1;
  ram[36110]  = 1;
  ram[36111]  = 1;
  ram[36112]  = 1;
  ram[36113]  = 0;
  ram[36114]  = 0;
  ram[36115]  = 1;
  ram[36116]  = 1;
  ram[36117]  = 1;
  ram[36118]  = 1;
  ram[36119]  = 1;
  ram[36120]  = 1;
  ram[36121]  = 1;
  ram[36122]  = 1;
  ram[36123]  = 1;
  ram[36124]  = 1;
  ram[36125]  = 1;
  ram[36126]  = 0;
  ram[36127]  = 0;
  ram[36128]  = 1;
  ram[36129]  = 1;
  ram[36130]  = 0;
  ram[36131]  = 1;
  ram[36132]  = 1;
  ram[36133]  = 1;
  ram[36134]  = 1;
  ram[36135]  = 1;
  ram[36136]  = 0;
  ram[36137]  = 1;
  ram[36138]  = 1;
  ram[36139]  = 0;
  ram[36140]  = 0;
  ram[36141]  = 1;
  ram[36142]  = 1;
  ram[36143]  = 1;
  ram[36144]  = 1;
  ram[36145]  = 1;
  ram[36146]  = 1;
  ram[36147]  = 0;
  ram[36148]  = 1;
  ram[36149]  = 1;
  ram[36150]  = 1;
  ram[36151]  = 0;
  ram[36152]  = 1;
  ram[36153]  = 0;
  ram[36154]  = 1;
  ram[36155]  = 1;
  ram[36156]  = 1;
  ram[36157]  = 0;
  ram[36158]  = 1;
  ram[36159]  = 0;
  ram[36160]  = 1;
  ram[36161]  = 1;
  ram[36162]  = 1;
  ram[36163]  = 1;
  ram[36164]  = 0;
  ram[36165]  = 1;
  ram[36166]  = 1;
  ram[36167]  = 1;
  ram[36168]  = 1;
  ram[36169]  = 1;
  ram[36170]  = 0;
  ram[36171]  = 1;
  ram[36172]  = 1;
  ram[36173]  = 1;
  ram[36174]  = 1;
  ram[36175]  = 1;
  ram[36176]  = 1;
  ram[36177]  = 1;
  ram[36178]  = 0;
  ram[36179]  = 0;
  ram[36180]  = 1;
  ram[36181]  = 1;
  ram[36182]  = 1;
  ram[36183]  = 1;
  ram[36184]  = 1;
  ram[36185]  = 1;
  ram[36186]  = 0;
  ram[36187]  = 1;
  ram[36188]  = 1;
  ram[36189]  = 1;
  ram[36190]  = 0;
  ram[36191]  = 1;
  ram[36192]  = 1;
  ram[36193]  = 1;
  ram[36194]  = 1;
  ram[36195]  = 1;
  ram[36196]  = 0;
  ram[36197]  = 1;
  ram[36198]  = 1;
  ram[36199]  = 1;
  ram[36200]  = 1;
  ram[36201]  = 1;
  ram[36202]  = 1;
  ram[36203]  = 1;
  ram[36204]  = 1;
  ram[36205]  = 0;
  ram[36206]  = 1;
  ram[36207]  = 1;
  ram[36208]  = 1;
  ram[36209]  = 1;
  ram[36210]  = 1;
  ram[36211]  = 0;
  ram[36212]  = 1;
  ram[36213]  = 1;
  ram[36214]  = 1;
  ram[36215]  = 1;
  ram[36216]  = 1;
  ram[36217]  = 0;
  ram[36218]  = 1;
  ram[36219]  = 1;
  ram[36220]  = 0;
  ram[36221]  = 0;
  ram[36222]  = 1;
  ram[36223]  = 1;
  ram[36224]  = 1;
  ram[36225]  = 1;
  ram[36226]  = 1;
  ram[36227]  = 1;
  ram[36228]  = 1;
  ram[36229]  = 1;
  ram[36230]  = 1;
  ram[36231]  = 1;
  ram[36232]  = 1;
  ram[36233]  = 1;
  ram[36234]  = 1;
  ram[36235]  = 0;
  ram[36236]  = 0;
  ram[36237]  = 1;
  ram[36238]  = 1;
  ram[36239]  = 1;
  ram[36240]  = 1;
  ram[36241]  = 1;
  ram[36242]  = 0;
  ram[36243]  = 0;
  ram[36244]  = 1;
  ram[36245]  = 1;
  ram[36246]  = 0;
  ram[36247]  = 1;
  ram[36248]  = 1;
  ram[36249]  = 1;
  ram[36250]  = 1;
  ram[36251]  = 1;
  ram[36252]  = 1;
  ram[36253]  = 0;
  ram[36254]  = 1;
  ram[36255]  = 1;
  ram[36256]  = 0;
  ram[36257]  = 0;
  ram[36258]  = 1;
  ram[36259]  = 1;
  ram[36260]  = 1;
  ram[36261]  = 1;
  ram[36262]  = 0;
  ram[36263]  = 1;
  ram[36264]  = 1;
  ram[36265]  = 1;
  ram[36266]  = 0;
  ram[36267]  = 1;
  ram[36268]  = 1;
  ram[36269]  = 1;
  ram[36270]  = 1;
  ram[36271]  = 1;
  ram[36272]  = 0;
  ram[36273]  = 1;
  ram[36274]  = 1;
  ram[36275]  = 1;
  ram[36276]  = 1;
  ram[36277]  = 1;
  ram[36278]  = 1;
  ram[36279]  = 0;
  ram[36280]  = 1;
  ram[36281]  = 1;
  ram[36282]  = 1;
  ram[36283]  = 1;
  ram[36284]  = 1;
  ram[36285]  = 1;
  ram[36286]  = 1;
  ram[36287]  = 1;
  ram[36288]  = 1;
  ram[36289]  = 1;
  ram[36290]  = 1;
  ram[36291]  = 1;
  ram[36292]  = 1;
  ram[36293]  = 1;
  ram[36294]  = 1;
  ram[36295]  = 1;
  ram[36296]  = 1;
  ram[36297]  = 1;
  ram[36298]  = 1;
  ram[36299]  = 1;
  ram[36300]  = 1;
  ram[36301]  = 1;
  ram[36302]  = 1;
  ram[36303]  = 1;
  ram[36304]  = 1;
  ram[36305]  = 1;
  ram[36306]  = 1;
  ram[36307]  = 1;
  ram[36308]  = 1;
  ram[36309]  = 1;
  ram[36310]  = 1;
  ram[36311]  = 1;
  ram[36312]  = 1;
  ram[36313]  = 1;
  ram[36314]  = 1;
  ram[36315]  = 1;
  ram[36316]  = 1;
  ram[36317]  = 0;
  ram[36318]  = 1;
  ram[36319]  = 1;
  ram[36320]  = 1;
  ram[36321]  = 1;
  ram[36322]  = 1;
  ram[36323]  = 0;
  ram[36324]  = 0;
  ram[36325]  = 1;
  ram[36326]  = 1;
  ram[36327]  = 1;
  ram[36328]  = 1;
  ram[36329]  = 1;
  ram[36330]  = 1;
  ram[36331]  = 0;
  ram[36332]  = 1;
  ram[36333]  = 1;
  ram[36334]  = 0;
  ram[36335]  = 0;
  ram[36336]  = 1;
  ram[36337]  = 1;
  ram[36338]  = 1;
  ram[36339]  = 1;
  ram[36340]  = 0;
  ram[36341]  = 0;
  ram[36342]  = 1;
  ram[36343]  = 1;
  ram[36344]  = 1;
  ram[36345]  = 0;
  ram[36346]  = 1;
  ram[36347]  = 1;
  ram[36348]  = 1;
  ram[36349]  = 1;
  ram[36350]  = 1;
  ram[36351]  = 1;
  ram[36352]  = 1;
  ram[36353]  = 1;
  ram[36354]  = 1;
  ram[36355]  = 1;
  ram[36356]  = 1;
  ram[36357]  = 1;
  ram[36358]  = 1;
  ram[36359]  = 1;
  ram[36360]  = 1;
  ram[36361]  = 1;
  ram[36362]  = 0;
  ram[36363]  = 1;
  ram[36364]  = 1;
  ram[36365]  = 0;
  ram[36366]  = 1;
  ram[36367]  = 1;
  ram[36368]  = 1;
  ram[36369]  = 1;
  ram[36370]  = 1;
  ram[36371]  = 1;
  ram[36372]  = 1;
  ram[36373]  = 1;
  ram[36374]  = 0;
  ram[36375]  = 1;
  ram[36376]  = 1;
  ram[36377]  = 1;
  ram[36378]  = 1;
  ram[36379]  = 1;
  ram[36380]  = 1;
  ram[36381]  = 0;
  ram[36382]  = 1;
  ram[36383]  = 1;
  ram[36384]  = 1;
  ram[36385]  = 0;
  ram[36386]  = 1;
  ram[36387]  = 1;
  ram[36388]  = 1;
  ram[36389]  = 1;
  ram[36390]  = 0;
  ram[36391]  = 0;
  ram[36392]  = 1;
  ram[36393]  = 1;
  ram[36394]  = 1;
  ram[36395]  = 1;
  ram[36396]  = 1;
  ram[36397]  = 1;
  ram[36398]  = 1;
  ram[36399]  = 1;
  ram[36400]  = 1;
  ram[36401]  = 1;
  ram[36402]  = 1;
  ram[36403]  = 1;
  ram[36404]  = 1;
  ram[36405]  = 0;
  ram[36406]  = 0;
  ram[36407]  = 1;
  ram[36408]  = 1;
  ram[36409]  = 1;
  ram[36410]  = 1;
  ram[36411]  = 1;
  ram[36412]  = 1;
  ram[36413]  = 1;
  ram[36414]  = 0;
  ram[36415]  = 1;
  ram[36416]  = 1;
  ram[36417]  = 1;
  ram[36418]  = 1;
  ram[36419]  = 1;
  ram[36420]  = 1;
  ram[36421]  = 1;
  ram[36422]  = 1;
  ram[36423]  = 1;
  ram[36424]  = 1;
  ram[36425]  = 1;
  ram[36426]  = 0;
  ram[36427]  = 0;
  ram[36428]  = 1;
  ram[36429]  = 1;
  ram[36430]  = 0;
  ram[36431]  = 1;
  ram[36432]  = 1;
  ram[36433]  = 1;
  ram[36434]  = 1;
  ram[36435]  = 1;
  ram[36436]  = 0;
  ram[36437]  = 1;
  ram[36438]  = 1;
  ram[36439]  = 1;
  ram[36440]  = 0;
  ram[36441]  = 1;
  ram[36442]  = 1;
  ram[36443]  = 1;
  ram[36444]  = 1;
  ram[36445]  = 1;
  ram[36446]  = 1;
  ram[36447]  = 0;
  ram[36448]  = 1;
  ram[36449]  = 1;
  ram[36450]  = 1;
  ram[36451]  = 0;
  ram[36452]  = 1;
  ram[36453]  = 0;
  ram[36454]  = 1;
  ram[36455]  = 1;
  ram[36456]  = 1;
  ram[36457]  = 0;
  ram[36458]  = 1;
  ram[36459]  = 0;
  ram[36460]  = 1;
  ram[36461]  = 1;
  ram[36462]  = 1;
  ram[36463]  = 1;
  ram[36464]  = 0;
  ram[36465]  = 1;
  ram[36466]  = 1;
  ram[36467]  = 1;
  ram[36468]  = 1;
  ram[36469]  = 1;
  ram[36470]  = 0;
  ram[36471]  = 1;
  ram[36472]  = 1;
  ram[36473]  = 1;
  ram[36474]  = 1;
  ram[36475]  = 1;
  ram[36476]  = 1;
  ram[36477]  = 1;
  ram[36478]  = 0;
  ram[36479]  = 0;
  ram[36480]  = 1;
  ram[36481]  = 1;
  ram[36482]  = 1;
  ram[36483]  = 1;
  ram[36484]  = 1;
  ram[36485]  = 1;
  ram[36486]  = 0;
  ram[36487]  = 1;
  ram[36488]  = 1;
  ram[36489]  = 1;
  ram[36490]  = 0;
  ram[36491]  = 1;
  ram[36492]  = 1;
  ram[36493]  = 1;
  ram[36494]  = 1;
  ram[36495]  = 1;
  ram[36496]  = 0;
  ram[36497]  = 1;
  ram[36498]  = 1;
  ram[36499]  = 1;
  ram[36500]  = 1;
  ram[36501]  = 1;
  ram[36502]  = 1;
  ram[36503]  = 1;
  ram[36504]  = 1;
  ram[36505]  = 0;
  ram[36506]  = 1;
  ram[36507]  = 1;
  ram[36508]  = 1;
  ram[36509]  = 1;
  ram[36510]  = 1;
  ram[36511]  = 0;
  ram[36512]  = 1;
  ram[36513]  = 1;
  ram[36514]  = 1;
  ram[36515]  = 1;
  ram[36516]  = 1;
  ram[36517]  = 0;
  ram[36518]  = 1;
  ram[36519]  = 1;
  ram[36520]  = 0;
  ram[36521]  = 0;
  ram[36522]  = 1;
  ram[36523]  = 1;
  ram[36524]  = 1;
  ram[36525]  = 1;
  ram[36526]  = 1;
  ram[36527]  = 1;
  ram[36528]  = 1;
  ram[36529]  = 1;
  ram[36530]  = 1;
  ram[36531]  = 1;
  ram[36532]  = 1;
  ram[36533]  = 1;
  ram[36534]  = 1;
  ram[36535]  = 0;
  ram[36536]  = 0;
  ram[36537]  = 1;
  ram[36538]  = 1;
  ram[36539]  = 1;
  ram[36540]  = 1;
  ram[36541]  = 1;
  ram[36542]  = 0;
  ram[36543]  = 0;
  ram[36544]  = 1;
  ram[36545]  = 1;
  ram[36546]  = 0;
  ram[36547]  = 1;
  ram[36548]  = 1;
  ram[36549]  = 1;
  ram[36550]  = 1;
  ram[36551]  = 1;
  ram[36552]  = 1;
  ram[36553]  = 0;
  ram[36554]  = 1;
  ram[36555]  = 1;
  ram[36556]  = 0;
  ram[36557]  = 1;
  ram[36558]  = 1;
  ram[36559]  = 1;
  ram[36560]  = 1;
  ram[36561]  = 1;
  ram[36562]  = 0;
  ram[36563]  = 1;
  ram[36564]  = 1;
  ram[36565]  = 1;
  ram[36566]  = 0;
  ram[36567]  = 1;
  ram[36568]  = 1;
  ram[36569]  = 1;
  ram[36570]  = 1;
  ram[36571]  = 1;
  ram[36572]  = 0;
  ram[36573]  = 1;
  ram[36574]  = 1;
  ram[36575]  = 1;
  ram[36576]  = 1;
  ram[36577]  = 1;
  ram[36578]  = 1;
  ram[36579]  = 0;
  ram[36580]  = 1;
  ram[36581]  = 1;
  ram[36582]  = 1;
  ram[36583]  = 1;
  ram[36584]  = 1;
  ram[36585]  = 1;
  ram[36586]  = 1;
  ram[36587]  = 1;
  ram[36588]  = 1;
  ram[36589]  = 1;
  ram[36590]  = 1;
  ram[36591]  = 1;
  ram[36592]  = 1;
  ram[36593]  = 1;
  ram[36594]  = 1;
  ram[36595]  = 1;
  ram[36596]  = 1;
  ram[36597]  = 1;
  ram[36598]  = 1;
  ram[36599]  = 1;
  ram[36600]  = 1;
  ram[36601]  = 1;
  ram[36602]  = 1;
  ram[36603]  = 1;
  ram[36604]  = 1;
  ram[36605]  = 1;
  ram[36606]  = 1;
  ram[36607]  = 1;
  ram[36608]  = 1;
  ram[36609]  = 1;
  ram[36610]  = 1;
  ram[36611]  = 1;
  ram[36612]  = 1;
  ram[36613]  = 1;
  ram[36614]  = 1;
  ram[36615]  = 1;
  ram[36616]  = 1;
  ram[36617]  = 0;
  ram[36618]  = 1;
  ram[36619]  = 1;
  ram[36620]  = 1;
  ram[36621]  = 1;
  ram[36622]  = 1;
  ram[36623]  = 1;
  ram[36624]  = 0;
  ram[36625]  = 1;
  ram[36626]  = 1;
  ram[36627]  = 1;
  ram[36628]  = 1;
  ram[36629]  = 1;
  ram[36630]  = 1;
  ram[36631]  = 0;
  ram[36632]  = 1;
  ram[36633]  = 1;
  ram[36634]  = 0;
  ram[36635]  = 0;
  ram[36636]  = 1;
  ram[36637]  = 1;
  ram[36638]  = 1;
  ram[36639]  = 1;
  ram[36640]  = 0;
  ram[36641]  = 0;
  ram[36642]  = 1;
  ram[36643]  = 1;
  ram[36644]  = 1;
  ram[36645]  = 0;
  ram[36646]  = 1;
  ram[36647]  = 1;
  ram[36648]  = 1;
  ram[36649]  = 1;
  ram[36650]  = 1;
  ram[36651]  = 1;
  ram[36652]  = 1;
  ram[36653]  = 1;
  ram[36654]  = 1;
  ram[36655]  = 0;
  ram[36656]  = 0;
  ram[36657]  = 1;
  ram[36658]  = 1;
  ram[36659]  = 1;
  ram[36660]  = 1;
  ram[36661]  = 1;
  ram[36662]  = 0;
  ram[36663]  = 1;
  ram[36664]  = 1;
  ram[36665]  = 0;
  ram[36666]  = 1;
  ram[36667]  = 1;
  ram[36668]  = 1;
  ram[36669]  = 1;
  ram[36670]  = 1;
  ram[36671]  = 1;
  ram[36672]  = 1;
  ram[36673]  = 1;
  ram[36674]  = 0;
  ram[36675]  = 1;
  ram[36676]  = 1;
  ram[36677]  = 1;
  ram[36678]  = 1;
  ram[36679]  = 1;
  ram[36680]  = 1;
  ram[36681]  = 0;
  ram[36682]  = 1;
  ram[36683]  = 1;
  ram[36684]  = 1;
  ram[36685]  = 0;
  ram[36686]  = 1;
  ram[36687]  = 1;
  ram[36688]  = 1;
  ram[36689]  = 1;
  ram[36690]  = 1;
  ram[36691]  = 0;
  ram[36692]  = 1;
  ram[36693]  = 1;
  ram[36694]  = 1;
  ram[36695]  = 1;
  ram[36696]  = 1;
  ram[36697]  = 1;
  ram[36698]  = 1;
  ram[36699]  = 1;
  ram[36700]  = 1;
  ram[36701]  = 1;
  ram[36702]  = 1;
  ram[36703]  = 1;
  ram[36704]  = 1;
  ram[36705]  = 0;
  ram[36706]  = 0;
  ram[36707]  = 1;
  ram[36708]  = 1;
  ram[36709]  = 1;
  ram[36710]  = 1;
  ram[36711]  = 1;
  ram[36712]  = 1;
  ram[36713]  = 1;
  ram[36714]  = 0;
  ram[36715]  = 1;
  ram[36716]  = 1;
  ram[36717]  = 1;
  ram[36718]  = 1;
  ram[36719]  = 1;
  ram[36720]  = 1;
  ram[36721]  = 1;
  ram[36722]  = 1;
  ram[36723]  = 1;
  ram[36724]  = 1;
  ram[36725]  = 1;
  ram[36726]  = 1;
  ram[36727]  = 0;
  ram[36728]  = 1;
  ram[36729]  = 1;
  ram[36730]  = 0;
  ram[36731]  = 1;
  ram[36732]  = 1;
  ram[36733]  = 1;
  ram[36734]  = 1;
  ram[36735]  = 1;
  ram[36736]  = 0;
  ram[36737]  = 1;
  ram[36738]  = 1;
  ram[36739]  = 1;
  ram[36740]  = 0;
  ram[36741]  = 1;
  ram[36742]  = 1;
  ram[36743]  = 1;
  ram[36744]  = 1;
  ram[36745]  = 1;
  ram[36746]  = 1;
  ram[36747]  = 0;
  ram[36748]  = 1;
  ram[36749]  = 1;
  ram[36750]  = 1;
  ram[36751]  = 0;
  ram[36752]  = 1;
  ram[36753]  = 0;
  ram[36754]  = 1;
  ram[36755]  = 1;
  ram[36756]  = 1;
  ram[36757]  = 0;
  ram[36758]  = 1;
  ram[36759]  = 0;
  ram[36760]  = 1;
  ram[36761]  = 1;
  ram[36762]  = 1;
  ram[36763]  = 1;
  ram[36764]  = 0;
  ram[36765]  = 1;
  ram[36766]  = 1;
  ram[36767]  = 1;
  ram[36768]  = 1;
  ram[36769]  = 1;
  ram[36770]  = 0;
  ram[36771]  = 1;
  ram[36772]  = 1;
  ram[36773]  = 1;
  ram[36774]  = 1;
  ram[36775]  = 1;
  ram[36776]  = 1;
  ram[36777]  = 1;
  ram[36778]  = 1;
  ram[36779]  = 0;
  ram[36780]  = 1;
  ram[36781]  = 1;
  ram[36782]  = 1;
  ram[36783]  = 1;
  ram[36784]  = 1;
  ram[36785]  = 1;
  ram[36786]  = 0;
  ram[36787]  = 1;
  ram[36788]  = 1;
  ram[36789]  = 1;
  ram[36790]  = 0;
  ram[36791]  = 1;
  ram[36792]  = 1;
  ram[36793]  = 1;
  ram[36794]  = 1;
  ram[36795]  = 1;
  ram[36796]  = 0;
  ram[36797]  = 1;
  ram[36798]  = 1;
  ram[36799]  = 1;
  ram[36800]  = 1;
  ram[36801]  = 1;
  ram[36802]  = 1;
  ram[36803]  = 1;
  ram[36804]  = 1;
  ram[36805]  = 0;
  ram[36806]  = 1;
  ram[36807]  = 1;
  ram[36808]  = 1;
  ram[36809]  = 1;
  ram[36810]  = 1;
  ram[36811]  = 0;
  ram[36812]  = 1;
  ram[36813]  = 1;
  ram[36814]  = 1;
  ram[36815]  = 1;
  ram[36816]  = 1;
  ram[36817]  = 0;
  ram[36818]  = 1;
  ram[36819]  = 1;
  ram[36820]  = 0;
  ram[36821]  = 0;
  ram[36822]  = 1;
  ram[36823]  = 1;
  ram[36824]  = 1;
  ram[36825]  = 1;
  ram[36826]  = 1;
  ram[36827]  = 1;
  ram[36828]  = 1;
  ram[36829]  = 1;
  ram[36830]  = 1;
  ram[36831]  = 1;
  ram[36832]  = 1;
  ram[36833]  = 1;
  ram[36834]  = 1;
  ram[36835]  = 0;
  ram[36836]  = 0;
  ram[36837]  = 1;
  ram[36838]  = 1;
  ram[36839]  = 1;
  ram[36840]  = 1;
  ram[36841]  = 1;
  ram[36842]  = 0;
  ram[36843]  = 0;
  ram[36844]  = 1;
  ram[36845]  = 1;
  ram[36846]  = 0;
  ram[36847]  = 1;
  ram[36848]  = 1;
  ram[36849]  = 1;
  ram[36850]  = 1;
  ram[36851]  = 1;
  ram[36852]  = 1;
  ram[36853]  = 0;
  ram[36854]  = 1;
  ram[36855]  = 1;
  ram[36856]  = 0;
  ram[36857]  = 1;
  ram[36858]  = 1;
  ram[36859]  = 1;
  ram[36860]  = 1;
  ram[36861]  = 1;
  ram[36862]  = 0;
  ram[36863]  = 1;
  ram[36864]  = 1;
  ram[36865]  = 1;
  ram[36866]  = 0;
  ram[36867]  = 1;
  ram[36868]  = 1;
  ram[36869]  = 1;
  ram[36870]  = 1;
  ram[36871]  = 1;
  ram[36872]  = 0;
  ram[36873]  = 1;
  ram[36874]  = 1;
  ram[36875]  = 1;
  ram[36876]  = 1;
  ram[36877]  = 1;
  ram[36878]  = 1;
  ram[36879]  = 0;
  ram[36880]  = 1;
  ram[36881]  = 1;
  ram[36882]  = 1;
  ram[36883]  = 1;
  ram[36884]  = 1;
  ram[36885]  = 1;
  ram[36886]  = 1;
  ram[36887]  = 1;
  ram[36888]  = 1;
  ram[36889]  = 1;
  ram[36890]  = 1;
  ram[36891]  = 1;
  ram[36892]  = 1;
  ram[36893]  = 1;
  ram[36894]  = 1;
  ram[36895]  = 1;
  ram[36896]  = 1;
  ram[36897]  = 1;
  ram[36898]  = 1;
  ram[36899]  = 1;
  ram[36900]  = 1;
  ram[36901]  = 1;
  ram[36902]  = 1;
  ram[36903]  = 1;
  ram[36904]  = 1;
  ram[36905]  = 1;
  ram[36906]  = 1;
  ram[36907]  = 1;
  ram[36908]  = 1;
  ram[36909]  = 1;
  ram[36910]  = 1;
  ram[36911]  = 1;
  ram[36912]  = 1;
  ram[36913]  = 1;
  ram[36914]  = 1;
  ram[36915]  = 1;
  ram[36916]  = 1;
  ram[36917]  = 0;
  ram[36918]  = 1;
  ram[36919]  = 1;
  ram[36920]  = 1;
  ram[36921]  = 1;
  ram[36922]  = 1;
  ram[36923]  = 1;
  ram[36924]  = 0;
  ram[36925]  = 1;
  ram[36926]  = 1;
  ram[36927]  = 1;
  ram[36928]  = 1;
  ram[36929]  = 1;
  ram[36930]  = 0;
  ram[36931]  = 0;
  ram[36932]  = 1;
  ram[36933]  = 1;
  ram[36934]  = 1;
  ram[36935]  = 0;
  ram[36936]  = 1;
  ram[36937]  = 1;
  ram[36938]  = 1;
  ram[36939]  = 1;
  ram[36940]  = 0;
  ram[36941]  = 0;
  ram[36942]  = 1;
  ram[36943]  = 1;
  ram[36944]  = 1;
  ram[36945]  = 0;
  ram[36946]  = 1;
  ram[36947]  = 1;
  ram[36948]  = 1;
  ram[36949]  = 1;
  ram[36950]  = 1;
  ram[36951]  = 1;
  ram[36952]  = 1;
  ram[36953]  = 1;
  ram[36954]  = 1;
  ram[36955]  = 1;
  ram[36956]  = 0;
  ram[36957]  = 1;
  ram[36958]  = 1;
  ram[36959]  = 1;
  ram[36960]  = 1;
  ram[36961]  = 1;
  ram[36962]  = 0;
  ram[36963]  = 1;
  ram[36964]  = 1;
  ram[36965]  = 0;
  ram[36966]  = 0;
  ram[36967]  = 1;
  ram[36968]  = 1;
  ram[36969]  = 1;
  ram[36970]  = 1;
  ram[36971]  = 0;
  ram[36972]  = 1;
  ram[36973]  = 1;
  ram[36974]  = 0;
  ram[36975]  = 1;
  ram[36976]  = 1;
  ram[36977]  = 1;
  ram[36978]  = 1;
  ram[36979]  = 1;
  ram[36980]  = 0;
  ram[36981]  = 0;
  ram[36982]  = 1;
  ram[36983]  = 1;
  ram[36984]  = 1;
  ram[36985]  = 0;
  ram[36986]  = 1;
  ram[36987]  = 1;
  ram[36988]  = 1;
  ram[36989]  = 1;
  ram[36990]  = 1;
  ram[36991]  = 0;
  ram[36992]  = 1;
  ram[36993]  = 1;
  ram[36994]  = 1;
  ram[36995]  = 1;
  ram[36996]  = 1;
  ram[36997]  = 0;
  ram[36998]  = 1;
  ram[36999]  = 1;
  ram[37000]  = 1;
  ram[37001]  = 1;
  ram[37002]  = 1;
  ram[37003]  = 1;
  ram[37004]  = 1;
  ram[37005]  = 0;
  ram[37006]  = 0;
  ram[37007]  = 1;
  ram[37008]  = 1;
  ram[37009]  = 0;
  ram[37010]  = 1;
  ram[37011]  = 1;
  ram[37012]  = 1;
  ram[37013]  = 1;
  ram[37014]  = 0;
  ram[37015]  = 1;
  ram[37016]  = 1;
  ram[37017]  = 1;
  ram[37018]  = 1;
  ram[37019]  = 1;
  ram[37020]  = 1;
  ram[37021]  = 0;
  ram[37022]  = 1;
  ram[37023]  = 1;
  ram[37024]  = 1;
  ram[37025]  = 1;
  ram[37026]  = 1;
  ram[37027]  = 0;
  ram[37028]  = 1;
  ram[37029]  = 1;
  ram[37030]  = 0;
  ram[37031]  = 1;
  ram[37032]  = 1;
  ram[37033]  = 1;
  ram[37034]  = 1;
  ram[37035]  = 1;
  ram[37036]  = 0;
  ram[37037]  = 1;
  ram[37038]  = 1;
  ram[37039]  = 1;
  ram[37040]  = 0;
  ram[37041]  = 1;
  ram[37042]  = 1;
  ram[37043]  = 1;
  ram[37044]  = 1;
  ram[37045]  = 1;
  ram[37046]  = 0;
  ram[37047]  = 0;
  ram[37048]  = 1;
  ram[37049]  = 1;
  ram[37050]  = 1;
  ram[37051]  = 0;
  ram[37052]  = 0;
  ram[37053]  = 0;
  ram[37054]  = 1;
  ram[37055]  = 1;
  ram[37056]  = 1;
  ram[37057]  = 0;
  ram[37058]  = 0;
  ram[37059]  = 0;
  ram[37060]  = 1;
  ram[37061]  = 1;
  ram[37062]  = 1;
  ram[37063]  = 1;
  ram[37064]  = 0;
  ram[37065]  = 1;
  ram[37066]  = 1;
  ram[37067]  = 1;
  ram[37068]  = 1;
  ram[37069]  = 1;
  ram[37070]  = 0;
  ram[37071]  = 1;
  ram[37072]  = 1;
  ram[37073]  = 1;
  ram[37074]  = 1;
  ram[37075]  = 1;
  ram[37076]  = 1;
  ram[37077]  = 1;
  ram[37078]  = 1;
  ram[37079]  = 0;
  ram[37080]  = 1;
  ram[37081]  = 1;
  ram[37082]  = 1;
  ram[37083]  = 1;
  ram[37084]  = 1;
  ram[37085]  = 0;
  ram[37086]  = 0;
  ram[37087]  = 1;
  ram[37088]  = 1;
  ram[37089]  = 1;
  ram[37090]  = 0;
  ram[37091]  = 1;
  ram[37092]  = 1;
  ram[37093]  = 1;
  ram[37094]  = 1;
  ram[37095]  = 1;
  ram[37096]  = 0;
  ram[37097]  = 1;
  ram[37098]  = 1;
  ram[37099]  = 1;
  ram[37100]  = 1;
  ram[37101]  = 1;
  ram[37102]  = 1;
  ram[37103]  = 1;
  ram[37104]  = 1;
  ram[37105]  = 0;
  ram[37106]  = 1;
  ram[37107]  = 1;
  ram[37108]  = 1;
  ram[37109]  = 1;
  ram[37110]  = 1;
  ram[37111]  = 0;
  ram[37112]  = 1;
  ram[37113]  = 1;
  ram[37114]  = 1;
  ram[37115]  = 1;
  ram[37116]  = 1;
  ram[37117]  = 0;
  ram[37118]  = 1;
  ram[37119]  = 1;
  ram[37120]  = 1;
  ram[37121]  = 0;
  ram[37122]  = 1;
  ram[37123]  = 1;
  ram[37124]  = 1;
  ram[37125]  = 1;
  ram[37126]  = 1;
  ram[37127]  = 0;
  ram[37128]  = 1;
  ram[37129]  = 1;
  ram[37130]  = 1;
  ram[37131]  = 1;
  ram[37132]  = 1;
  ram[37133]  = 1;
  ram[37134]  = 1;
  ram[37135]  = 1;
  ram[37136]  = 0;
  ram[37137]  = 1;
  ram[37138]  = 1;
  ram[37139]  = 1;
  ram[37140]  = 1;
  ram[37141]  = 1;
  ram[37142]  = 0;
  ram[37143]  = 1;
  ram[37144]  = 1;
  ram[37145]  = 1;
  ram[37146]  = 0;
  ram[37147]  = 1;
  ram[37148]  = 1;
  ram[37149]  = 1;
  ram[37150]  = 1;
  ram[37151]  = 1;
  ram[37152]  = 0;
  ram[37153]  = 0;
  ram[37154]  = 1;
  ram[37155]  = 1;
  ram[37156]  = 0;
  ram[37157]  = 1;
  ram[37158]  = 1;
  ram[37159]  = 1;
  ram[37160]  = 1;
  ram[37161]  = 0;
  ram[37162]  = 0;
  ram[37163]  = 1;
  ram[37164]  = 1;
  ram[37165]  = 1;
  ram[37166]  = 0;
  ram[37167]  = 1;
  ram[37168]  = 1;
  ram[37169]  = 1;
  ram[37170]  = 1;
  ram[37171]  = 1;
  ram[37172]  = 0;
  ram[37173]  = 0;
  ram[37174]  = 1;
  ram[37175]  = 1;
  ram[37176]  = 1;
  ram[37177]  = 1;
  ram[37178]  = 0;
  ram[37179]  = 0;
  ram[37180]  = 1;
  ram[37181]  = 1;
  ram[37182]  = 1;
  ram[37183]  = 1;
  ram[37184]  = 1;
  ram[37185]  = 1;
  ram[37186]  = 1;
  ram[37187]  = 1;
  ram[37188]  = 1;
  ram[37189]  = 1;
  ram[37190]  = 1;
  ram[37191]  = 1;
  ram[37192]  = 1;
  ram[37193]  = 1;
  ram[37194]  = 1;
  ram[37195]  = 1;
  ram[37196]  = 1;
  ram[37197]  = 1;
  ram[37198]  = 1;
  ram[37199]  = 1;
  ram[37200]  = 1;
  ram[37201]  = 1;
  ram[37202]  = 1;
  ram[37203]  = 1;
  ram[37204]  = 1;
  ram[37205]  = 1;
  ram[37206]  = 1;
  ram[37207]  = 1;
  ram[37208]  = 1;
  ram[37209]  = 1;
  ram[37210]  = 1;
  ram[37211]  = 1;
  ram[37212]  = 1;
  ram[37213]  = 1;
  ram[37214]  = 1;
  ram[37215]  = 1;
  ram[37216]  = 1;
  ram[37217]  = 0;
  ram[37218]  = 1;
  ram[37219]  = 1;
  ram[37220]  = 1;
  ram[37221]  = 1;
  ram[37222]  = 1;
  ram[37223]  = 1;
  ram[37224]  = 0;
  ram[37225]  = 0;
  ram[37226]  = 1;
  ram[37227]  = 1;
  ram[37228]  = 1;
  ram[37229]  = 1;
  ram[37230]  = 0;
  ram[37231]  = 1;
  ram[37232]  = 1;
  ram[37233]  = 1;
  ram[37234]  = 1;
  ram[37235]  = 0;
  ram[37236]  = 1;
  ram[37237]  = 1;
  ram[37238]  = 1;
  ram[37239]  = 1;
  ram[37240]  = 0;
  ram[37241]  = 0;
  ram[37242]  = 1;
  ram[37243]  = 1;
  ram[37244]  = 1;
  ram[37245]  = 0;
  ram[37246]  = 1;
  ram[37247]  = 1;
  ram[37248]  = 1;
  ram[37249]  = 1;
  ram[37250]  = 1;
  ram[37251]  = 1;
  ram[37252]  = 1;
  ram[37253]  = 1;
  ram[37254]  = 1;
  ram[37255]  = 1;
  ram[37256]  = 0;
  ram[37257]  = 1;
  ram[37258]  = 1;
  ram[37259]  = 1;
  ram[37260]  = 1;
  ram[37261]  = 0;
  ram[37262]  = 0;
  ram[37263]  = 1;
  ram[37264]  = 1;
  ram[37265]  = 1;
  ram[37266]  = 0;
  ram[37267]  = 1;
  ram[37268]  = 1;
  ram[37269]  = 1;
  ram[37270]  = 1;
  ram[37271]  = 0;
  ram[37272]  = 1;
  ram[37273]  = 1;
  ram[37274]  = 0;
  ram[37275]  = 0;
  ram[37276]  = 1;
  ram[37277]  = 1;
  ram[37278]  = 1;
  ram[37279]  = 1;
  ram[37280]  = 0;
  ram[37281]  = 1;
  ram[37282]  = 1;
  ram[37283]  = 1;
  ram[37284]  = 1;
  ram[37285]  = 0;
  ram[37286]  = 1;
  ram[37287]  = 1;
  ram[37288]  = 1;
  ram[37289]  = 1;
  ram[37290]  = 1;
  ram[37291]  = 0;
  ram[37292]  = 0;
  ram[37293]  = 1;
  ram[37294]  = 1;
  ram[37295]  = 1;
  ram[37296]  = 0;
  ram[37297]  = 0;
  ram[37298]  = 1;
  ram[37299]  = 1;
  ram[37300]  = 1;
  ram[37301]  = 1;
  ram[37302]  = 1;
  ram[37303]  = 1;
  ram[37304]  = 1;
  ram[37305]  = 0;
  ram[37306]  = 0;
  ram[37307]  = 1;
  ram[37308]  = 1;
  ram[37309]  = 0;
  ram[37310]  = 1;
  ram[37311]  = 1;
  ram[37312]  = 1;
  ram[37313]  = 1;
  ram[37314]  = 0;
  ram[37315]  = 1;
  ram[37316]  = 1;
  ram[37317]  = 1;
  ram[37318]  = 1;
  ram[37319]  = 1;
  ram[37320]  = 1;
  ram[37321]  = 0;
  ram[37322]  = 0;
  ram[37323]  = 1;
  ram[37324]  = 1;
  ram[37325]  = 1;
  ram[37326]  = 0;
  ram[37327]  = 0;
  ram[37328]  = 1;
  ram[37329]  = 1;
  ram[37330]  = 0;
  ram[37331]  = 1;
  ram[37332]  = 1;
  ram[37333]  = 1;
  ram[37334]  = 1;
  ram[37335]  = 1;
  ram[37336]  = 0;
  ram[37337]  = 1;
  ram[37338]  = 1;
  ram[37339]  = 1;
  ram[37340]  = 0;
  ram[37341]  = 0;
  ram[37342]  = 1;
  ram[37343]  = 1;
  ram[37344]  = 1;
  ram[37345]  = 1;
  ram[37346]  = 0;
  ram[37347]  = 1;
  ram[37348]  = 1;
  ram[37349]  = 1;
  ram[37350]  = 1;
  ram[37351]  = 1;
  ram[37352]  = 0;
  ram[37353]  = 0;
  ram[37354]  = 1;
  ram[37355]  = 1;
  ram[37356]  = 1;
  ram[37357]  = 0;
  ram[37358]  = 0;
  ram[37359]  = 1;
  ram[37360]  = 1;
  ram[37361]  = 1;
  ram[37362]  = 1;
  ram[37363]  = 1;
  ram[37364]  = 0;
  ram[37365]  = 1;
  ram[37366]  = 1;
  ram[37367]  = 1;
  ram[37368]  = 1;
  ram[37369]  = 1;
  ram[37370]  = 0;
  ram[37371]  = 1;
  ram[37372]  = 1;
  ram[37373]  = 1;
  ram[37374]  = 1;
  ram[37375]  = 1;
  ram[37376]  = 1;
  ram[37377]  = 1;
  ram[37378]  = 1;
  ram[37379]  = 0;
  ram[37380]  = 0;
  ram[37381]  = 1;
  ram[37382]  = 1;
  ram[37383]  = 1;
  ram[37384]  = 1;
  ram[37385]  = 0;
  ram[37386]  = 1;
  ram[37387]  = 1;
  ram[37388]  = 1;
  ram[37389]  = 1;
  ram[37390]  = 0;
  ram[37391]  = 1;
  ram[37392]  = 1;
  ram[37393]  = 1;
  ram[37394]  = 1;
  ram[37395]  = 1;
  ram[37396]  = 0;
  ram[37397]  = 1;
  ram[37398]  = 1;
  ram[37399]  = 1;
  ram[37400]  = 1;
  ram[37401]  = 1;
  ram[37402]  = 1;
  ram[37403]  = 1;
  ram[37404]  = 1;
  ram[37405]  = 0;
  ram[37406]  = 1;
  ram[37407]  = 1;
  ram[37408]  = 1;
  ram[37409]  = 1;
  ram[37410]  = 1;
  ram[37411]  = 0;
  ram[37412]  = 1;
  ram[37413]  = 1;
  ram[37414]  = 1;
  ram[37415]  = 1;
  ram[37416]  = 1;
  ram[37417]  = 0;
  ram[37418]  = 1;
  ram[37419]  = 1;
  ram[37420]  = 1;
  ram[37421]  = 0;
  ram[37422]  = 0;
  ram[37423]  = 1;
  ram[37424]  = 1;
  ram[37425]  = 1;
  ram[37426]  = 0;
  ram[37427]  = 0;
  ram[37428]  = 1;
  ram[37429]  = 1;
  ram[37430]  = 1;
  ram[37431]  = 1;
  ram[37432]  = 1;
  ram[37433]  = 1;
  ram[37434]  = 1;
  ram[37435]  = 0;
  ram[37436]  = 0;
  ram[37437]  = 0;
  ram[37438]  = 1;
  ram[37439]  = 1;
  ram[37440]  = 1;
  ram[37441]  = 1;
  ram[37442]  = 0;
  ram[37443]  = 1;
  ram[37444]  = 1;
  ram[37445]  = 1;
  ram[37446]  = 0;
  ram[37447]  = 0;
  ram[37448]  = 1;
  ram[37449]  = 1;
  ram[37450]  = 1;
  ram[37451]  = 1;
  ram[37452]  = 0;
  ram[37453]  = 0;
  ram[37454]  = 1;
  ram[37455]  = 1;
  ram[37456]  = 0;
  ram[37457]  = 0;
  ram[37458]  = 1;
  ram[37459]  = 1;
  ram[37460]  = 1;
  ram[37461]  = 0;
  ram[37462]  = 0;
  ram[37463]  = 1;
  ram[37464]  = 1;
  ram[37465]  = 1;
  ram[37466]  = 0;
  ram[37467]  = 1;
  ram[37468]  = 1;
  ram[37469]  = 1;
  ram[37470]  = 1;
  ram[37471]  = 1;
  ram[37472]  = 1;
  ram[37473]  = 0;
  ram[37474]  = 1;
  ram[37475]  = 1;
  ram[37476]  = 1;
  ram[37477]  = 1;
  ram[37478]  = 0;
  ram[37479]  = 0;
  ram[37480]  = 1;
  ram[37481]  = 1;
  ram[37482]  = 1;
  ram[37483]  = 1;
  ram[37484]  = 1;
  ram[37485]  = 1;
  ram[37486]  = 1;
  ram[37487]  = 1;
  ram[37488]  = 1;
  ram[37489]  = 1;
  ram[37490]  = 1;
  ram[37491]  = 1;
  ram[37492]  = 1;
  ram[37493]  = 1;
  ram[37494]  = 1;
  ram[37495]  = 1;
  ram[37496]  = 1;
  ram[37497]  = 1;
  ram[37498]  = 1;
  ram[37499]  = 1;
  ram[37500]  = 1;
  ram[37501]  = 1;
  ram[37502]  = 1;
  ram[37503]  = 1;
  ram[37504]  = 1;
  ram[37505]  = 1;
  ram[37506]  = 1;
  ram[37507]  = 1;
  ram[37508]  = 1;
  ram[37509]  = 1;
  ram[37510]  = 1;
  ram[37511]  = 1;
  ram[37512]  = 1;
  ram[37513]  = 1;
  ram[37514]  = 1;
  ram[37515]  = 1;
  ram[37516]  = 1;
  ram[37517]  = 0;
  ram[37518]  = 1;
  ram[37519]  = 1;
  ram[37520]  = 1;
  ram[37521]  = 1;
  ram[37522]  = 1;
  ram[37523]  = 1;
  ram[37524]  = 1;
  ram[37525]  = 0;
  ram[37526]  = 0;
  ram[37527]  = 1;
  ram[37528]  = 1;
  ram[37529]  = 0;
  ram[37530]  = 0;
  ram[37531]  = 1;
  ram[37532]  = 1;
  ram[37533]  = 1;
  ram[37534]  = 1;
  ram[37535]  = 0;
  ram[37536]  = 0;
  ram[37537]  = 1;
  ram[37538]  = 1;
  ram[37539]  = 0;
  ram[37540]  = 1;
  ram[37541]  = 0;
  ram[37542]  = 1;
  ram[37543]  = 1;
  ram[37544]  = 1;
  ram[37545]  = 0;
  ram[37546]  = 1;
  ram[37547]  = 1;
  ram[37548]  = 1;
  ram[37549]  = 1;
  ram[37550]  = 1;
  ram[37551]  = 1;
  ram[37552]  = 1;
  ram[37553]  = 1;
  ram[37554]  = 1;
  ram[37555]  = 1;
  ram[37556]  = 0;
  ram[37557]  = 0;
  ram[37558]  = 1;
  ram[37559]  = 1;
  ram[37560]  = 0;
  ram[37561]  = 0;
  ram[37562]  = 1;
  ram[37563]  = 1;
  ram[37564]  = 1;
  ram[37565]  = 1;
  ram[37566]  = 0;
  ram[37567]  = 0;
  ram[37568]  = 1;
  ram[37569]  = 1;
  ram[37570]  = 0;
  ram[37571]  = 0;
  ram[37572]  = 1;
  ram[37573]  = 1;
  ram[37574]  = 1;
  ram[37575]  = 0;
  ram[37576]  = 0;
  ram[37577]  = 1;
  ram[37578]  = 1;
  ram[37579]  = 0;
  ram[37580]  = 0;
  ram[37581]  = 1;
  ram[37582]  = 1;
  ram[37583]  = 1;
  ram[37584]  = 1;
  ram[37585]  = 0;
  ram[37586]  = 1;
  ram[37587]  = 1;
  ram[37588]  = 1;
  ram[37589]  = 1;
  ram[37590]  = 1;
  ram[37591]  = 1;
  ram[37592]  = 0;
  ram[37593]  = 0;
  ram[37594]  = 1;
  ram[37595]  = 0;
  ram[37596]  = 0;
  ram[37597]  = 1;
  ram[37598]  = 1;
  ram[37599]  = 1;
  ram[37600]  = 1;
  ram[37601]  = 1;
  ram[37602]  = 1;
  ram[37603]  = 1;
  ram[37604]  = 1;
  ram[37605]  = 0;
  ram[37606]  = 0;
  ram[37607]  = 1;
  ram[37608]  = 1;
  ram[37609]  = 0;
  ram[37610]  = 0;
  ram[37611]  = 1;
  ram[37612]  = 1;
  ram[37613]  = 0;
  ram[37614]  = 0;
  ram[37615]  = 1;
  ram[37616]  = 1;
  ram[37617]  = 1;
  ram[37618]  = 1;
  ram[37619]  = 1;
  ram[37620]  = 1;
  ram[37621]  = 1;
  ram[37622]  = 0;
  ram[37623]  = 1;
  ram[37624]  = 1;
  ram[37625]  = 1;
  ram[37626]  = 0;
  ram[37627]  = 1;
  ram[37628]  = 1;
  ram[37629]  = 1;
  ram[37630]  = 0;
  ram[37631]  = 1;
  ram[37632]  = 1;
  ram[37633]  = 1;
  ram[37634]  = 1;
  ram[37635]  = 1;
  ram[37636]  = 0;
  ram[37637]  = 1;
  ram[37638]  = 1;
  ram[37639]  = 1;
  ram[37640]  = 1;
  ram[37641]  = 0;
  ram[37642]  = 0;
  ram[37643]  = 1;
  ram[37644]  = 1;
  ram[37645]  = 0;
  ram[37646]  = 0;
  ram[37647]  = 1;
  ram[37648]  = 1;
  ram[37649]  = 1;
  ram[37650]  = 1;
  ram[37651]  = 1;
  ram[37652]  = 0;
  ram[37653]  = 1;
  ram[37654]  = 1;
  ram[37655]  = 1;
  ram[37656]  = 1;
  ram[37657]  = 1;
  ram[37658]  = 0;
  ram[37659]  = 1;
  ram[37660]  = 1;
  ram[37661]  = 1;
  ram[37662]  = 1;
  ram[37663]  = 1;
  ram[37664]  = 0;
  ram[37665]  = 1;
  ram[37666]  = 1;
  ram[37667]  = 1;
  ram[37668]  = 1;
  ram[37669]  = 1;
  ram[37670]  = 0;
  ram[37671]  = 1;
  ram[37672]  = 1;
  ram[37673]  = 1;
  ram[37674]  = 1;
  ram[37675]  = 1;
  ram[37676]  = 1;
  ram[37677]  = 1;
  ram[37678]  = 1;
  ram[37679]  = 1;
  ram[37680]  = 0;
  ram[37681]  = 0;
  ram[37682]  = 1;
  ram[37683]  = 1;
  ram[37684]  = 0;
  ram[37685]  = 0;
  ram[37686]  = 1;
  ram[37687]  = 1;
  ram[37688]  = 1;
  ram[37689]  = 1;
  ram[37690]  = 0;
  ram[37691]  = 1;
  ram[37692]  = 1;
  ram[37693]  = 1;
  ram[37694]  = 1;
  ram[37695]  = 1;
  ram[37696]  = 0;
  ram[37697]  = 1;
  ram[37698]  = 1;
  ram[37699]  = 1;
  ram[37700]  = 1;
  ram[37701]  = 1;
  ram[37702]  = 1;
  ram[37703]  = 1;
  ram[37704]  = 1;
  ram[37705]  = 0;
  ram[37706]  = 0;
  ram[37707]  = 1;
  ram[37708]  = 1;
  ram[37709]  = 1;
  ram[37710]  = 1;
  ram[37711]  = 0;
  ram[37712]  = 1;
  ram[37713]  = 1;
  ram[37714]  = 1;
  ram[37715]  = 1;
  ram[37716]  = 1;
  ram[37717]  = 0;
  ram[37718]  = 1;
  ram[37719]  = 1;
  ram[37720]  = 1;
  ram[37721]  = 1;
  ram[37722]  = 0;
  ram[37723]  = 0;
  ram[37724]  = 1;
  ram[37725]  = 0;
  ram[37726]  = 0;
  ram[37727]  = 1;
  ram[37728]  = 1;
  ram[37729]  = 1;
  ram[37730]  = 1;
  ram[37731]  = 1;
  ram[37732]  = 1;
  ram[37733]  = 1;
  ram[37734]  = 1;
  ram[37735]  = 0;
  ram[37736]  = 0;
  ram[37737]  = 0;
  ram[37738]  = 0;
  ram[37739]  = 1;
  ram[37740]  = 0;
  ram[37741]  = 0;
  ram[37742]  = 1;
  ram[37743]  = 1;
  ram[37744]  = 1;
  ram[37745]  = 1;
  ram[37746]  = 1;
  ram[37747]  = 0;
  ram[37748]  = 0;
  ram[37749]  = 1;
  ram[37750]  = 1;
  ram[37751]  = 0;
  ram[37752]  = 0;
  ram[37753]  = 1;
  ram[37754]  = 1;
  ram[37755]  = 1;
  ram[37756]  = 1;
  ram[37757]  = 0;
  ram[37758]  = 1;
  ram[37759]  = 1;
  ram[37760]  = 0;
  ram[37761]  = 1;
  ram[37762]  = 0;
  ram[37763]  = 1;
  ram[37764]  = 1;
  ram[37765]  = 1;
  ram[37766]  = 0;
  ram[37767]  = 1;
  ram[37768]  = 1;
  ram[37769]  = 1;
  ram[37770]  = 1;
  ram[37771]  = 1;
  ram[37772]  = 1;
  ram[37773]  = 0;
  ram[37774]  = 0;
  ram[37775]  = 1;
  ram[37776]  = 1;
  ram[37777]  = 0;
  ram[37778]  = 1;
  ram[37779]  = 0;
  ram[37780]  = 1;
  ram[37781]  = 1;
  ram[37782]  = 1;
  ram[37783]  = 1;
  ram[37784]  = 1;
  ram[37785]  = 1;
  ram[37786]  = 1;
  ram[37787]  = 1;
  ram[37788]  = 1;
  ram[37789]  = 1;
  ram[37790]  = 1;
  ram[37791]  = 1;
  ram[37792]  = 1;
  ram[37793]  = 1;
  ram[37794]  = 1;
  ram[37795]  = 1;
  ram[37796]  = 1;
  ram[37797]  = 1;
  ram[37798]  = 1;
  ram[37799]  = 1;
  ram[37800]  = 1;
  ram[37801]  = 1;
  ram[37802]  = 1;
  ram[37803]  = 1;
  ram[37804]  = 1;
  ram[37805]  = 1;
  ram[37806]  = 1;
  ram[37807]  = 1;
  ram[37808]  = 1;
  ram[37809]  = 1;
  ram[37810]  = 1;
  ram[37811]  = 1;
  ram[37812]  = 1;
  ram[37813]  = 1;
  ram[37814]  = 1;
  ram[37815]  = 1;
  ram[37816]  = 1;
  ram[37817]  = 0;
  ram[37818]  = 1;
  ram[37819]  = 1;
  ram[37820]  = 1;
  ram[37821]  = 1;
  ram[37822]  = 1;
  ram[37823]  = 1;
  ram[37824]  = 1;
  ram[37825]  = 1;
  ram[37826]  = 0;
  ram[37827]  = 0;
  ram[37828]  = 0;
  ram[37829]  = 0;
  ram[37830]  = 1;
  ram[37831]  = 1;
  ram[37832]  = 1;
  ram[37833]  = 1;
  ram[37834]  = 1;
  ram[37835]  = 1;
  ram[37836]  = 0;
  ram[37837]  = 0;
  ram[37838]  = 0;
  ram[37839]  = 1;
  ram[37840]  = 1;
  ram[37841]  = 0;
  ram[37842]  = 1;
  ram[37843]  = 1;
  ram[37844]  = 1;
  ram[37845]  = 0;
  ram[37846]  = 1;
  ram[37847]  = 1;
  ram[37848]  = 1;
  ram[37849]  = 1;
  ram[37850]  = 1;
  ram[37851]  = 1;
  ram[37852]  = 1;
  ram[37853]  = 1;
  ram[37854]  = 1;
  ram[37855]  = 1;
  ram[37856]  = 1;
  ram[37857]  = 0;
  ram[37858]  = 0;
  ram[37859]  = 0;
  ram[37860]  = 0;
  ram[37861]  = 0;
  ram[37862]  = 1;
  ram[37863]  = 1;
  ram[37864]  = 1;
  ram[37865]  = 1;
  ram[37866]  = 1;
  ram[37867]  = 0;
  ram[37868]  = 0;
  ram[37869]  = 0;
  ram[37870]  = 0;
  ram[37871]  = 1;
  ram[37872]  = 1;
  ram[37873]  = 1;
  ram[37874]  = 1;
  ram[37875]  = 1;
  ram[37876]  = 0;
  ram[37877]  = 0;
  ram[37878]  = 0;
  ram[37879]  = 0;
  ram[37880]  = 1;
  ram[37881]  = 1;
  ram[37882]  = 1;
  ram[37883]  = 1;
  ram[37884]  = 1;
  ram[37885]  = 0;
  ram[37886]  = 1;
  ram[37887]  = 1;
  ram[37888]  = 1;
  ram[37889]  = 1;
  ram[37890]  = 1;
  ram[37891]  = 1;
  ram[37892]  = 0;
  ram[37893]  = 0;
  ram[37894]  = 0;
  ram[37895]  = 0;
  ram[37896]  = 0;
  ram[37897]  = 1;
  ram[37898]  = 1;
  ram[37899]  = 1;
  ram[37900]  = 1;
  ram[37901]  = 1;
  ram[37902]  = 1;
  ram[37903]  = 1;
  ram[37904]  = 1;
  ram[37905]  = 0;
  ram[37906]  = 0;
  ram[37907]  = 1;
  ram[37908]  = 1;
  ram[37909]  = 1;
  ram[37910]  = 0;
  ram[37911]  = 0;
  ram[37912]  = 0;
  ram[37913]  = 0;
  ram[37914]  = 1;
  ram[37915]  = 1;
  ram[37916]  = 1;
  ram[37917]  = 1;
  ram[37918]  = 1;
  ram[37919]  = 1;
  ram[37920]  = 1;
  ram[37921]  = 1;
  ram[37922]  = 0;
  ram[37923]  = 0;
  ram[37924]  = 0;
  ram[37925]  = 0;
  ram[37926]  = 0;
  ram[37927]  = 1;
  ram[37928]  = 1;
  ram[37929]  = 1;
  ram[37930]  = 0;
  ram[37931]  = 1;
  ram[37932]  = 1;
  ram[37933]  = 1;
  ram[37934]  = 1;
  ram[37935]  = 1;
  ram[37936]  = 0;
  ram[37937]  = 1;
  ram[37938]  = 1;
  ram[37939]  = 1;
  ram[37940]  = 1;
  ram[37941]  = 1;
  ram[37942]  = 0;
  ram[37943]  = 0;
  ram[37944]  = 0;
  ram[37945]  = 0;
  ram[37946]  = 1;
  ram[37947]  = 1;
  ram[37948]  = 1;
  ram[37949]  = 1;
  ram[37950]  = 1;
  ram[37951]  = 1;
  ram[37952]  = 0;
  ram[37953]  = 1;
  ram[37954]  = 1;
  ram[37955]  = 1;
  ram[37956]  = 1;
  ram[37957]  = 1;
  ram[37958]  = 0;
  ram[37959]  = 1;
  ram[37960]  = 1;
  ram[37961]  = 1;
  ram[37962]  = 1;
  ram[37963]  = 1;
  ram[37964]  = 0;
  ram[37965]  = 1;
  ram[37966]  = 1;
  ram[37967]  = 1;
  ram[37968]  = 1;
  ram[37969]  = 1;
  ram[37970]  = 0;
  ram[37971]  = 1;
  ram[37972]  = 1;
  ram[37973]  = 1;
  ram[37974]  = 1;
  ram[37975]  = 1;
  ram[37976]  = 1;
  ram[37977]  = 1;
  ram[37978]  = 1;
  ram[37979]  = 1;
  ram[37980]  = 0;
  ram[37981]  = 0;
  ram[37982]  = 0;
  ram[37983]  = 0;
  ram[37984]  = 0;
  ram[37985]  = 1;
  ram[37986]  = 1;
  ram[37987]  = 1;
  ram[37988]  = 1;
  ram[37989]  = 0;
  ram[37990]  = 0;
  ram[37991]  = 1;
  ram[37992]  = 1;
  ram[37993]  = 1;
  ram[37994]  = 1;
  ram[37995]  = 1;
  ram[37996]  = 0;
  ram[37997]  = 1;
  ram[37998]  = 1;
  ram[37999]  = 1;
  ram[38000]  = 1;
  ram[38001]  = 1;
  ram[38002]  = 1;
  ram[38003]  = 1;
  ram[38004]  = 1;
  ram[38005]  = 1;
  ram[38006]  = 0;
  ram[38007]  = 0;
  ram[38008]  = 0;
  ram[38009]  = 1;
  ram[38010]  = 1;
  ram[38011]  = 0;
  ram[38012]  = 1;
  ram[38013]  = 1;
  ram[38014]  = 1;
  ram[38015]  = 1;
  ram[38016]  = 1;
  ram[38017]  = 0;
  ram[38018]  = 1;
  ram[38019]  = 1;
  ram[38020]  = 1;
  ram[38021]  = 1;
  ram[38022]  = 0;
  ram[38023]  = 0;
  ram[38024]  = 0;
  ram[38025]  = 0;
  ram[38026]  = 1;
  ram[38027]  = 1;
  ram[38028]  = 1;
  ram[38029]  = 1;
  ram[38030]  = 1;
  ram[38031]  = 1;
  ram[38032]  = 1;
  ram[38033]  = 1;
  ram[38034]  = 1;
  ram[38035]  = 0;
  ram[38036]  = 0;
  ram[38037]  = 1;
  ram[38038]  = 0;
  ram[38039]  = 0;
  ram[38040]  = 0;
  ram[38041]  = 0;
  ram[38042]  = 1;
  ram[38043]  = 1;
  ram[38044]  = 1;
  ram[38045]  = 1;
  ram[38046]  = 1;
  ram[38047]  = 1;
  ram[38048]  = 0;
  ram[38049]  = 0;
  ram[38050]  = 0;
  ram[38051]  = 0;
  ram[38052]  = 1;
  ram[38053]  = 1;
  ram[38054]  = 1;
  ram[38055]  = 1;
  ram[38056]  = 1;
  ram[38057]  = 0;
  ram[38058]  = 0;
  ram[38059]  = 0;
  ram[38060]  = 0;
  ram[38061]  = 1;
  ram[38062]  = 0;
  ram[38063]  = 1;
  ram[38064]  = 1;
  ram[38065]  = 1;
  ram[38066]  = 0;
  ram[38067]  = 1;
  ram[38068]  = 1;
  ram[38069]  = 1;
  ram[38070]  = 1;
  ram[38071]  = 1;
  ram[38072]  = 1;
  ram[38073]  = 1;
  ram[38074]  = 0;
  ram[38075]  = 0;
  ram[38076]  = 0;
  ram[38077]  = 0;
  ram[38078]  = 1;
  ram[38079]  = 0;
  ram[38080]  = 1;
  ram[38081]  = 1;
  ram[38082]  = 1;
  ram[38083]  = 1;
  ram[38084]  = 1;
  ram[38085]  = 1;
  ram[38086]  = 1;
  ram[38087]  = 1;
  ram[38088]  = 1;
  ram[38089]  = 1;
  ram[38090]  = 1;
  ram[38091]  = 1;
  ram[38092]  = 1;
  ram[38093]  = 1;
  ram[38094]  = 1;
  ram[38095]  = 1;
  ram[38096]  = 1;
  ram[38097]  = 1;
  ram[38098]  = 1;
  ram[38099]  = 1;
  ram[38100]  = 1;
  ram[38101]  = 1;
  ram[38102]  = 1;
  ram[38103]  = 1;
  ram[38104]  = 1;
  ram[38105]  = 1;
  ram[38106]  = 1;
  ram[38107]  = 1;
  ram[38108]  = 1;
  ram[38109]  = 1;
  ram[38110]  = 1;
  ram[38111]  = 1;
  ram[38112]  = 1;
  ram[38113]  = 1;
  ram[38114]  = 1;
  ram[38115]  = 1;
  ram[38116]  = 1;
  ram[38117]  = 1;
  ram[38118]  = 1;
  ram[38119]  = 1;
  ram[38120]  = 1;
  ram[38121]  = 1;
  ram[38122]  = 1;
  ram[38123]  = 1;
  ram[38124]  = 1;
  ram[38125]  = 1;
  ram[38126]  = 1;
  ram[38127]  = 1;
  ram[38128]  = 1;
  ram[38129]  = 1;
  ram[38130]  = 1;
  ram[38131]  = 1;
  ram[38132]  = 1;
  ram[38133]  = 1;
  ram[38134]  = 1;
  ram[38135]  = 1;
  ram[38136]  = 1;
  ram[38137]  = 1;
  ram[38138]  = 1;
  ram[38139]  = 1;
  ram[38140]  = 1;
  ram[38141]  = 1;
  ram[38142]  = 1;
  ram[38143]  = 1;
  ram[38144]  = 1;
  ram[38145]  = 1;
  ram[38146]  = 1;
  ram[38147]  = 1;
  ram[38148]  = 1;
  ram[38149]  = 1;
  ram[38150]  = 1;
  ram[38151]  = 1;
  ram[38152]  = 1;
  ram[38153]  = 1;
  ram[38154]  = 1;
  ram[38155]  = 1;
  ram[38156]  = 1;
  ram[38157]  = 1;
  ram[38158]  = 1;
  ram[38159]  = 1;
  ram[38160]  = 1;
  ram[38161]  = 1;
  ram[38162]  = 1;
  ram[38163]  = 1;
  ram[38164]  = 1;
  ram[38165]  = 1;
  ram[38166]  = 1;
  ram[38167]  = 1;
  ram[38168]  = 1;
  ram[38169]  = 1;
  ram[38170]  = 1;
  ram[38171]  = 1;
  ram[38172]  = 1;
  ram[38173]  = 1;
  ram[38174]  = 1;
  ram[38175]  = 1;
  ram[38176]  = 1;
  ram[38177]  = 1;
  ram[38178]  = 1;
  ram[38179]  = 1;
  ram[38180]  = 1;
  ram[38181]  = 1;
  ram[38182]  = 1;
  ram[38183]  = 1;
  ram[38184]  = 1;
  ram[38185]  = 1;
  ram[38186]  = 1;
  ram[38187]  = 1;
  ram[38188]  = 1;
  ram[38189]  = 1;
  ram[38190]  = 1;
  ram[38191]  = 1;
  ram[38192]  = 1;
  ram[38193]  = 1;
  ram[38194]  = 1;
  ram[38195]  = 1;
  ram[38196]  = 1;
  ram[38197]  = 1;
  ram[38198]  = 1;
  ram[38199]  = 1;
  ram[38200]  = 1;
  ram[38201]  = 1;
  ram[38202]  = 1;
  ram[38203]  = 1;
  ram[38204]  = 1;
  ram[38205]  = 1;
  ram[38206]  = 1;
  ram[38207]  = 1;
  ram[38208]  = 1;
  ram[38209]  = 1;
  ram[38210]  = 1;
  ram[38211]  = 1;
  ram[38212]  = 1;
  ram[38213]  = 1;
  ram[38214]  = 1;
  ram[38215]  = 1;
  ram[38216]  = 1;
  ram[38217]  = 1;
  ram[38218]  = 1;
  ram[38219]  = 1;
  ram[38220]  = 1;
  ram[38221]  = 1;
  ram[38222]  = 1;
  ram[38223]  = 1;
  ram[38224]  = 1;
  ram[38225]  = 1;
  ram[38226]  = 1;
  ram[38227]  = 1;
  ram[38228]  = 1;
  ram[38229]  = 1;
  ram[38230]  = 1;
  ram[38231]  = 1;
  ram[38232]  = 1;
  ram[38233]  = 1;
  ram[38234]  = 1;
  ram[38235]  = 1;
  ram[38236]  = 1;
  ram[38237]  = 1;
  ram[38238]  = 1;
  ram[38239]  = 1;
  ram[38240]  = 1;
  ram[38241]  = 1;
  ram[38242]  = 1;
  ram[38243]  = 1;
  ram[38244]  = 1;
  ram[38245]  = 1;
  ram[38246]  = 1;
  ram[38247]  = 1;
  ram[38248]  = 1;
  ram[38249]  = 1;
  ram[38250]  = 1;
  ram[38251]  = 1;
  ram[38252]  = 1;
  ram[38253]  = 1;
  ram[38254]  = 1;
  ram[38255]  = 1;
  ram[38256]  = 1;
  ram[38257]  = 1;
  ram[38258]  = 1;
  ram[38259]  = 1;
  ram[38260]  = 1;
  ram[38261]  = 1;
  ram[38262]  = 1;
  ram[38263]  = 1;
  ram[38264]  = 1;
  ram[38265]  = 1;
  ram[38266]  = 1;
  ram[38267]  = 1;
  ram[38268]  = 1;
  ram[38269]  = 1;
  ram[38270]  = 1;
  ram[38271]  = 1;
  ram[38272]  = 1;
  ram[38273]  = 1;
  ram[38274]  = 1;
  ram[38275]  = 1;
  ram[38276]  = 1;
  ram[38277]  = 1;
  ram[38278]  = 1;
  ram[38279]  = 1;
  ram[38280]  = 1;
  ram[38281]  = 1;
  ram[38282]  = 1;
  ram[38283]  = 1;
  ram[38284]  = 1;
  ram[38285]  = 1;
  ram[38286]  = 1;
  ram[38287]  = 1;
  ram[38288]  = 1;
  ram[38289]  = 1;
  ram[38290]  = 1;
  ram[38291]  = 1;
  ram[38292]  = 1;
  ram[38293]  = 1;
  ram[38294]  = 1;
  ram[38295]  = 1;
  ram[38296]  = 1;
  ram[38297]  = 1;
  ram[38298]  = 1;
  ram[38299]  = 1;
  ram[38300]  = 1;
  ram[38301]  = 1;
  ram[38302]  = 1;
  ram[38303]  = 1;
  ram[38304]  = 1;
  ram[38305]  = 1;
  ram[38306]  = 1;
  ram[38307]  = 1;
  ram[38308]  = 1;
  ram[38309]  = 1;
  ram[38310]  = 1;
  ram[38311]  = 1;
  ram[38312]  = 1;
  ram[38313]  = 1;
  ram[38314]  = 1;
  ram[38315]  = 1;
  ram[38316]  = 1;
  ram[38317]  = 1;
  ram[38318]  = 1;
  ram[38319]  = 1;
  ram[38320]  = 1;
  ram[38321]  = 1;
  ram[38322]  = 1;
  ram[38323]  = 1;
  ram[38324]  = 1;
  ram[38325]  = 1;
  ram[38326]  = 1;
  ram[38327]  = 1;
  ram[38328]  = 1;
  ram[38329]  = 1;
  ram[38330]  = 1;
  ram[38331]  = 1;
  ram[38332]  = 1;
  ram[38333]  = 1;
  ram[38334]  = 1;
  ram[38335]  = 1;
  ram[38336]  = 1;
  ram[38337]  = 1;
  ram[38338]  = 1;
  ram[38339]  = 1;
  ram[38340]  = 1;
  ram[38341]  = 1;
  ram[38342]  = 1;
  ram[38343]  = 1;
  ram[38344]  = 1;
  ram[38345]  = 1;
  ram[38346]  = 1;
  ram[38347]  = 1;
  ram[38348]  = 1;
  ram[38349]  = 1;
  ram[38350]  = 1;
  ram[38351]  = 1;
  ram[38352]  = 1;
  ram[38353]  = 1;
  ram[38354]  = 1;
  ram[38355]  = 1;
  ram[38356]  = 1;
  ram[38357]  = 1;
  ram[38358]  = 1;
  ram[38359]  = 1;
  ram[38360]  = 1;
  ram[38361]  = 1;
  ram[38362]  = 1;
  ram[38363]  = 1;
  ram[38364]  = 1;
  ram[38365]  = 1;
  ram[38366]  = 1;
  ram[38367]  = 1;
  ram[38368]  = 1;
  ram[38369]  = 1;
  ram[38370]  = 1;
  ram[38371]  = 1;
  ram[38372]  = 1;
  ram[38373]  = 1;
  ram[38374]  = 1;
  ram[38375]  = 1;
  ram[38376]  = 1;
  ram[38377]  = 1;
  ram[38378]  = 1;
  ram[38379]  = 1;
  ram[38380]  = 1;
  ram[38381]  = 1;
  ram[38382]  = 1;
  ram[38383]  = 1;
  ram[38384]  = 1;
  ram[38385]  = 1;
  ram[38386]  = 1;
  ram[38387]  = 1;
  ram[38388]  = 1;
  ram[38389]  = 1;
  ram[38390]  = 1;
  ram[38391]  = 1;
  ram[38392]  = 1;
  ram[38393]  = 1;
  ram[38394]  = 1;
  ram[38395]  = 1;
  ram[38396]  = 1;
  ram[38397]  = 1;
  ram[38398]  = 1;
  ram[38399]  = 1;
  ram[38400]  = 1;
  ram[38401]  = 1;
  ram[38402]  = 1;
  ram[38403]  = 1;
  ram[38404]  = 1;
  ram[38405]  = 1;
  ram[38406]  = 1;
  ram[38407]  = 1;
  ram[38408]  = 1;
  ram[38409]  = 1;
  ram[38410]  = 1;
  ram[38411]  = 1;
  ram[38412]  = 1;
  ram[38413]  = 1;
  ram[38414]  = 1;
  ram[38415]  = 1;
  ram[38416]  = 1;
  ram[38417]  = 1;
  ram[38418]  = 1;
  ram[38419]  = 1;
  ram[38420]  = 1;
  ram[38421]  = 1;
  ram[38422]  = 1;
  ram[38423]  = 1;
  ram[38424]  = 1;
  ram[38425]  = 1;
  ram[38426]  = 1;
  ram[38427]  = 1;
  ram[38428]  = 1;
  ram[38429]  = 1;
  ram[38430]  = 1;
  ram[38431]  = 1;
  ram[38432]  = 1;
  ram[38433]  = 1;
  ram[38434]  = 1;
  ram[38435]  = 1;
  ram[38436]  = 1;
  ram[38437]  = 1;
  ram[38438]  = 1;
  ram[38439]  = 1;
  ram[38440]  = 1;
  ram[38441]  = 1;
  ram[38442]  = 1;
  ram[38443]  = 1;
  ram[38444]  = 1;
  ram[38445]  = 1;
  ram[38446]  = 1;
  ram[38447]  = 1;
  ram[38448]  = 1;
  ram[38449]  = 1;
  ram[38450]  = 1;
  ram[38451]  = 1;
  ram[38452]  = 1;
  ram[38453]  = 1;
  ram[38454]  = 1;
  ram[38455]  = 1;
  ram[38456]  = 1;
  ram[38457]  = 1;
  ram[38458]  = 1;
  ram[38459]  = 1;
  ram[38460]  = 1;
  ram[38461]  = 1;
  ram[38462]  = 1;
  ram[38463]  = 1;
  ram[38464]  = 1;
  ram[38465]  = 1;
  ram[38466]  = 1;
  ram[38467]  = 1;
  ram[38468]  = 1;
  ram[38469]  = 1;
  ram[38470]  = 1;
  ram[38471]  = 1;
  ram[38472]  = 1;
  ram[38473]  = 1;
  ram[38474]  = 1;
  ram[38475]  = 1;
  ram[38476]  = 1;
  ram[38477]  = 1;
  ram[38478]  = 1;
  ram[38479]  = 1;
  ram[38480]  = 1;
  ram[38481]  = 1;
  ram[38482]  = 1;
  ram[38483]  = 1;
  ram[38484]  = 1;
  ram[38485]  = 1;
  ram[38486]  = 1;
  ram[38487]  = 1;
  ram[38488]  = 1;
  ram[38489]  = 1;
  ram[38490]  = 1;
  ram[38491]  = 1;
  ram[38492]  = 1;
  ram[38493]  = 1;
  ram[38494]  = 1;
  ram[38495]  = 1;
  ram[38496]  = 1;
  ram[38497]  = 1;
  ram[38498]  = 1;
  ram[38499]  = 1;
  ram[38500]  = 1;
  ram[38501]  = 1;
  ram[38502]  = 1;
  ram[38503]  = 1;
  ram[38504]  = 1;
  ram[38505]  = 1;
  ram[38506]  = 1;
  ram[38507]  = 1;
  ram[38508]  = 1;
  ram[38509]  = 1;
  ram[38510]  = 1;
  ram[38511]  = 1;
  ram[38512]  = 1;
  ram[38513]  = 1;
  ram[38514]  = 1;
  ram[38515]  = 1;
  ram[38516]  = 1;
  ram[38517]  = 1;
  ram[38518]  = 1;
  ram[38519]  = 1;
  ram[38520]  = 1;
  ram[38521]  = 1;
  ram[38522]  = 1;
  ram[38523]  = 1;
  ram[38524]  = 1;
  ram[38525]  = 1;
  ram[38526]  = 1;
  ram[38527]  = 1;
  ram[38528]  = 1;
  ram[38529]  = 1;
  ram[38530]  = 1;
  ram[38531]  = 1;
  ram[38532]  = 1;
  ram[38533]  = 1;
  ram[38534]  = 1;
  ram[38535]  = 1;
  ram[38536]  = 1;
  ram[38537]  = 1;
  ram[38538]  = 1;
  ram[38539]  = 1;
  ram[38540]  = 1;
  ram[38541]  = 1;
  ram[38542]  = 1;
  ram[38543]  = 1;
  ram[38544]  = 1;
  ram[38545]  = 1;
  ram[38546]  = 1;
  ram[38547]  = 1;
  ram[38548]  = 1;
  ram[38549]  = 1;
  ram[38550]  = 1;
  ram[38551]  = 1;
  ram[38552]  = 1;
  ram[38553]  = 1;
  ram[38554]  = 1;
  ram[38555]  = 1;
  ram[38556]  = 1;
  ram[38557]  = 1;
  ram[38558]  = 1;
  ram[38559]  = 1;
  ram[38560]  = 1;
  ram[38561]  = 1;
  ram[38562]  = 1;
  ram[38563]  = 1;
  ram[38564]  = 1;
  ram[38565]  = 1;
  ram[38566]  = 1;
  ram[38567]  = 1;
  ram[38568]  = 1;
  ram[38569]  = 1;
  ram[38570]  = 1;
  ram[38571]  = 1;
  ram[38572]  = 1;
  ram[38573]  = 1;
  ram[38574]  = 1;
  ram[38575]  = 1;
  ram[38576]  = 1;
  ram[38577]  = 1;
  ram[38578]  = 1;
  ram[38579]  = 1;
  ram[38580]  = 1;
  ram[38581]  = 1;
  ram[38582]  = 1;
  ram[38583]  = 1;
  ram[38584]  = 1;
  ram[38585]  = 1;
  ram[38586]  = 1;
  ram[38587]  = 1;
  ram[38588]  = 1;
  ram[38589]  = 1;
  ram[38590]  = 1;
  ram[38591]  = 1;
  ram[38592]  = 1;
  ram[38593]  = 1;
  ram[38594]  = 1;
  ram[38595]  = 1;
  ram[38596]  = 1;
  ram[38597]  = 1;
  ram[38598]  = 1;
  ram[38599]  = 1;
  ram[38600]  = 1;
  ram[38601]  = 1;
  ram[38602]  = 1;
  ram[38603]  = 1;
  ram[38604]  = 1;
  ram[38605]  = 1;
  ram[38606]  = 1;
  ram[38607]  = 1;
  ram[38608]  = 1;
  ram[38609]  = 1;
  ram[38610]  = 1;
  ram[38611]  = 1;
  ram[38612]  = 1;
  ram[38613]  = 1;
  ram[38614]  = 1;
  ram[38615]  = 1;
  ram[38616]  = 1;
  ram[38617]  = 1;
  ram[38618]  = 1;
  ram[38619]  = 1;
  ram[38620]  = 1;
  ram[38621]  = 1;
  ram[38622]  = 1;
  ram[38623]  = 1;
  ram[38624]  = 1;
  ram[38625]  = 1;
  ram[38626]  = 1;
  ram[38627]  = 1;
  ram[38628]  = 1;
  ram[38629]  = 1;
  ram[38630]  = 1;
  ram[38631]  = 1;
  ram[38632]  = 1;
  ram[38633]  = 1;
  ram[38634]  = 1;
  ram[38635]  = 1;
  ram[38636]  = 1;
  ram[38637]  = 1;
  ram[38638]  = 1;
  ram[38639]  = 1;
  ram[38640]  = 1;
  ram[38641]  = 1;
  ram[38642]  = 1;
  ram[38643]  = 1;
  ram[38644]  = 1;
  ram[38645]  = 1;
  ram[38646]  = 1;
  ram[38647]  = 1;
  ram[38648]  = 1;
  ram[38649]  = 1;
  ram[38650]  = 1;
  ram[38651]  = 1;
  ram[38652]  = 1;
  ram[38653]  = 1;
  ram[38654]  = 1;
  ram[38655]  = 1;
  ram[38656]  = 1;
  ram[38657]  = 1;
  ram[38658]  = 1;
  ram[38659]  = 1;
  ram[38660]  = 1;
  ram[38661]  = 1;
  ram[38662]  = 1;
  ram[38663]  = 1;
  ram[38664]  = 1;
  ram[38665]  = 1;
  ram[38666]  = 1;
  ram[38667]  = 1;
  ram[38668]  = 1;
  ram[38669]  = 1;
  ram[38670]  = 1;
  ram[38671]  = 1;
  ram[38672]  = 1;
  ram[38673]  = 1;
  ram[38674]  = 1;
  ram[38675]  = 1;
  ram[38676]  = 1;
  ram[38677]  = 1;
  ram[38678]  = 1;
  ram[38679]  = 1;
  ram[38680]  = 1;
  ram[38681]  = 1;
  ram[38682]  = 1;
  ram[38683]  = 1;
  ram[38684]  = 1;
  ram[38685]  = 1;
  ram[38686]  = 1;
  ram[38687]  = 1;
  ram[38688]  = 1;
  ram[38689]  = 1;
  ram[38690]  = 1;
  ram[38691]  = 1;
  ram[38692]  = 1;
  ram[38693]  = 1;
  ram[38694]  = 1;
  ram[38695]  = 1;
  ram[38696]  = 1;
  ram[38697]  = 1;
  ram[38698]  = 1;
  ram[38699]  = 1;
  ram[38700]  = 1;
  ram[38701]  = 1;
  ram[38702]  = 1;
  ram[38703]  = 1;
  ram[38704]  = 1;
  ram[38705]  = 1;
  ram[38706]  = 1;
  ram[38707]  = 1;
  ram[38708]  = 1;
  ram[38709]  = 1;
  ram[38710]  = 1;
  ram[38711]  = 1;
  ram[38712]  = 1;
  ram[38713]  = 1;
  ram[38714]  = 1;
  ram[38715]  = 1;
  ram[38716]  = 1;
  ram[38717]  = 1;
  ram[38718]  = 1;
  ram[38719]  = 1;
  ram[38720]  = 1;
  ram[38721]  = 1;
  ram[38722]  = 1;
  ram[38723]  = 1;
  ram[38724]  = 1;
  ram[38725]  = 1;
  ram[38726]  = 1;
  ram[38727]  = 1;
  ram[38728]  = 1;
  ram[38729]  = 1;
  ram[38730]  = 1;
  ram[38731]  = 1;
  ram[38732]  = 1;
  ram[38733]  = 1;
  ram[38734]  = 1;
  ram[38735]  = 1;
  ram[38736]  = 1;
  ram[38737]  = 1;
  ram[38738]  = 1;
  ram[38739]  = 1;
  ram[38740]  = 1;
  ram[38741]  = 1;
  ram[38742]  = 1;
  ram[38743]  = 1;
  ram[38744]  = 1;
  ram[38745]  = 1;
  ram[38746]  = 1;
  ram[38747]  = 1;
  ram[38748]  = 1;
  ram[38749]  = 1;
  ram[38750]  = 1;
  ram[38751]  = 1;
  ram[38752]  = 1;
  ram[38753]  = 1;
  ram[38754]  = 1;
  ram[38755]  = 1;
  ram[38756]  = 1;
  ram[38757]  = 1;
  ram[38758]  = 1;
  ram[38759]  = 1;
  ram[38760]  = 1;
  ram[38761]  = 1;
  ram[38762]  = 1;
  ram[38763]  = 1;
  ram[38764]  = 1;
  ram[38765]  = 1;
  ram[38766]  = 1;
  ram[38767]  = 1;
  ram[38768]  = 1;
  ram[38769]  = 1;
  ram[38770]  = 1;
  ram[38771]  = 1;
  ram[38772]  = 1;
  ram[38773]  = 1;
  ram[38774]  = 1;
  ram[38775]  = 1;
  ram[38776]  = 1;
  ram[38777]  = 1;
  ram[38778]  = 1;
  ram[38779]  = 1;
  ram[38780]  = 1;
  ram[38781]  = 1;
  ram[38782]  = 1;
  ram[38783]  = 1;
  ram[38784]  = 1;
  ram[38785]  = 1;
  ram[38786]  = 1;
  ram[38787]  = 1;
  ram[38788]  = 1;
  ram[38789]  = 1;
  ram[38790]  = 1;
  ram[38791]  = 1;
  ram[38792]  = 1;
  ram[38793]  = 1;
  ram[38794]  = 1;
  ram[38795]  = 1;
  ram[38796]  = 1;
  ram[38797]  = 1;
  ram[38798]  = 1;
  ram[38799]  = 1;
  ram[38800]  = 1;
  ram[38801]  = 1;
  ram[38802]  = 1;
  ram[38803]  = 1;
  ram[38804]  = 1;
  ram[38805]  = 1;
  ram[38806]  = 1;
  ram[38807]  = 1;
  ram[38808]  = 1;
  ram[38809]  = 1;
  ram[38810]  = 1;
  ram[38811]  = 1;
  ram[38812]  = 1;
  ram[38813]  = 1;
  ram[38814]  = 1;
  ram[38815]  = 1;
  ram[38816]  = 1;
  ram[38817]  = 1;
  ram[38818]  = 1;
  ram[38819]  = 1;
  ram[38820]  = 1;
  ram[38821]  = 1;
  ram[38822]  = 1;
  ram[38823]  = 1;
  ram[38824]  = 1;
  ram[38825]  = 1;
  ram[38826]  = 1;
  ram[38827]  = 1;
  ram[38828]  = 1;
  ram[38829]  = 1;
  ram[38830]  = 1;
  ram[38831]  = 1;
  ram[38832]  = 1;
  ram[38833]  = 1;
  ram[38834]  = 1;
  ram[38835]  = 1;
  ram[38836]  = 1;
  ram[38837]  = 1;
  ram[38838]  = 1;
  ram[38839]  = 1;
  ram[38840]  = 1;
  ram[38841]  = 1;
  ram[38842]  = 1;
  ram[38843]  = 1;
  ram[38844]  = 1;
  ram[38845]  = 1;
  ram[38846]  = 1;
  ram[38847]  = 1;
  ram[38848]  = 1;
  ram[38849]  = 1;
  ram[38850]  = 1;
  ram[38851]  = 1;
  ram[38852]  = 1;
  ram[38853]  = 1;
  ram[38854]  = 1;
  ram[38855]  = 1;
  ram[38856]  = 1;
  ram[38857]  = 1;
  ram[38858]  = 1;
  ram[38859]  = 1;
  ram[38860]  = 1;
  ram[38861]  = 1;
  ram[38862]  = 1;
  ram[38863]  = 1;
  ram[38864]  = 1;
  ram[38865]  = 1;
  ram[38866]  = 1;
  ram[38867]  = 1;
  ram[38868]  = 1;
  ram[38869]  = 1;
  ram[38870]  = 1;
  ram[38871]  = 1;
  ram[38872]  = 1;
  ram[38873]  = 1;
  ram[38874]  = 1;
  ram[38875]  = 1;
  ram[38876]  = 1;
  ram[38877]  = 1;
  ram[38878]  = 1;
  ram[38879]  = 1;
  ram[38880]  = 1;
  ram[38881]  = 1;
  ram[38882]  = 1;
  ram[38883]  = 1;
  ram[38884]  = 1;
  ram[38885]  = 1;
  ram[38886]  = 1;
  ram[38887]  = 1;
  ram[38888]  = 1;
  ram[38889]  = 1;
  ram[38890]  = 1;
  ram[38891]  = 1;
  ram[38892]  = 1;
  ram[38893]  = 1;
  ram[38894]  = 1;
  ram[38895]  = 1;
  ram[38896]  = 1;
  ram[38897]  = 1;
  ram[38898]  = 1;
  ram[38899]  = 1;
  ram[38900]  = 1;
  ram[38901]  = 1;
  ram[38902]  = 1;
  ram[38903]  = 1;
  ram[38904]  = 1;
  ram[38905]  = 1;
  ram[38906]  = 1;
  ram[38907]  = 1;
  ram[38908]  = 1;
  ram[38909]  = 1;
  ram[38910]  = 1;
  ram[38911]  = 1;
  ram[38912]  = 1;
  ram[38913]  = 1;
  ram[38914]  = 1;
  ram[38915]  = 1;
  ram[38916]  = 1;
  ram[38917]  = 1;
  ram[38918]  = 1;
  ram[38919]  = 1;
  ram[38920]  = 1;
  ram[38921]  = 1;
  ram[38922]  = 1;
  ram[38923]  = 1;
  ram[38924]  = 1;
  ram[38925]  = 1;
  ram[38926]  = 1;
  ram[38927]  = 1;
  ram[38928]  = 1;
  ram[38929]  = 1;
  ram[38930]  = 1;
  ram[38931]  = 1;
  ram[38932]  = 1;
  ram[38933]  = 1;
  ram[38934]  = 1;
  ram[38935]  = 1;
  ram[38936]  = 1;
  ram[38937]  = 1;
  ram[38938]  = 1;
  ram[38939]  = 1;
  ram[38940]  = 1;
  ram[38941]  = 1;
  ram[38942]  = 1;
  ram[38943]  = 1;
  ram[38944]  = 1;
  ram[38945]  = 1;
  ram[38946]  = 1;
  ram[38947]  = 1;
  ram[38948]  = 1;
  ram[38949]  = 1;
  ram[38950]  = 1;
  ram[38951]  = 1;
  ram[38952]  = 1;
  ram[38953]  = 1;
  ram[38954]  = 1;
  ram[38955]  = 1;
  ram[38956]  = 1;
  ram[38957]  = 1;
  ram[38958]  = 1;
  ram[38959]  = 1;
  ram[38960]  = 1;
  ram[38961]  = 1;
  ram[38962]  = 1;
  ram[38963]  = 1;
  ram[38964]  = 1;
  ram[38965]  = 1;
  ram[38966]  = 1;
  ram[38967]  = 1;
  ram[38968]  = 1;
  ram[38969]  = 1;
  ram[38970]  = 1;
  ram[38971]  = 1;
  ram[38972]  = 1;
  ram[38973]  = 1;
  ram[38974]  = 1;
  ram[38975]  = 1;
  ram[38976]  = 1;
  ram[38977]  = 1;
  ram[38978]  = 1;
  ram[38979]  = 1;
  ram[38980]  = 1;
  ram[38981]  = 1;
  ram[38982]  = 1;
  ram[38983]  = 1;
  ram[38984]  = 1;
  ram[38985]  = 1;
  ram[38986]  = 1;
  ram[38987]  = 1;
  ram[38988]  = 1;
  ram[38989]  = 1;
  ram[38990]  = 1;
  ram[38991]  = 1;
  ram[38992]  = 1;
  ram[38993]  = 1;
  ram[38994]  = 1;
  ram[38995]  = 1;
  ram[38996]  = 1;
  ram[38997]  = 1;
  ram[38998]  = 1;
  ram[38999]  = 1;
  ram[39000]  = 1;
  ram[39001]  = 1;
  ram[39002]  = 1;
  ram[39003]  = 1;
  ram[39004]  = 1;
  ram[39005]  = 1;
  ram[39006]  = 1;
  ram[39007]  = 1;
  ram[39008]  = 1;
  ram[39009]  = 1;
  ram[39010]  = 1;
  ram[39011]  = 1;
  ram[39012]  = 1;
  ram[39013]  = 1;
  ram[39014]  = 1;
  ram[39015]  = 1;
  ram[39016]  = 1;
  ram[39017]  = 1;
  ram[39018]  = 1;
  ram[39019]  = 1;
  ram[39020]  = 1;
  ram[39021]  = 1;
  ram[39022]  = 1;
  ram[39023]  = 1;
  ram[39024]  = 1;
  ram[39025]  = 1;
  ram[39026]  = 1;
  ram[39027]  = 1;
  ram[39028]  = 1;
  ram[39029]  = 1;
  ram[39030]  = 1;
  ram[39031]  = 1;
  ram[39032]  = 1;
  ram[39033]  = 1;
  ram[39034]  = 1;
  ram[39035]  = 1;
  ram[39036]  = 1;
  ram[39037]  = 1;
  ram[39038]  = 1;
  ram[39039]  = 1;
  ram[39040]  = 1;
  ram[39041]  = 1;
  ram[39042]  = 1;
  ram[39043]  = 1;
  ram[39044]  = 1;
  ram[39045]  = 1;
  ram[39046]  = 1;
  ram[39047]  = 1;
  ram[39048]  = 1;
  ram[39049]  = 1;
  ram[39050]  = 1;
  ram[39051]  = 1;
  ram[39052]  = 1;
  ram[39053]  = 1;
  ram[39054]  = 1;
  ram[39055]  = 1;
  ram[39056]  = 1;
  ram[39057]  = 1;
  ram[39058]  = 1;
  ram[39059]  = 1;
  ram[39060]  = 1;
  ram[39061]  = 1;
  ram[39062]  = 1;
  ram[39063]  = 1;
  ram[39064]  = 1;
  ram[39065]  = 1;
  ram[39066]  = 1;
  ram[39067]  = 1;
  ram[39068]  = 1;
  ram[39069]  = 1;
  ram[39070]  = 1;
  ram[39071]  = 1;
  ram[39072]  = 1;
  ram[39073]  = 1;
  ram[39074]  = 1;
  ram[39075]  = 1;
  ram[39076]  = 1;
  ram[39077]  = 1;
  ram[39078]  = 1;
  ram[39079]  = 1;
  ram[39080]  = 1;
  ram[39081]  = 1;
  ram[39082]  = 1;
  ram[39083]  = 1;
  ram[39084]  = 1;
  ram[39085]  = 1;
  ram[39086]  = 1;
  ram[39087]  = 1;
  ram[39088]  = 1;
  ram[39089]  = 1;
  ram[39090]  = 1;
  ram[39091]  = 1;
  ram[39092]  = 1;
  ram[39093]  = 1;
  ram[39094]  = 1;
  ram[39095]  = 1;
  ram[39096]  = 1;
  ram[39097]  = 1;
  ram[39098]  = 1;
  ram[39099]  = 1;
  ram[39100]  = 1;
  ram[39101]  = 1;
  ram[39102]  = 1;
  ram[39103]  = 1;
  ram[39104]  = 1;
  ram[39105]  = 1;
  ram[39106]  = 1;
  ram[39107]  = 1;
  ram[39108]  = 1;
  ram[39109]  = 1;
  ram[39110]  = 1;
  ram[39111]  = 1;
  ram[39112]  = 1;
  ram[39113]  = 1;
  ram[39114]  = 1;
  ram[39115]  = 1;
  ram[39116]  = 1;
  ram[39117]  = 1;
  ram[39118]  = 1;
  ram[39119]  = 1;
  ram[39120]  = 1;
  ram[39121]  = 1;
  ram[39122]  = 1;
  ram[39123]  = 1;
  ram[39124]  = 1;
  ram[39125]  = 1;
  ram[39126]  = 1;
  ram[39127]  = 1;
  ram[39128]  = 1;
  ram[39129]  = 1;
  ram[39130]  = 1;
  ram[39131]  = 1;
  ram[39132]  = 1;
  ram[39133]  = 1;
  ram[39134]  = 1;
  ram[39135]  = 1;
  ram[39136]  = 1;
  ram[39137]  = 1;
  ram[39138]  = 1;
  ram[39139]  = 1;
  ram[39140]  = 1;
  ram[39141]  = 1;
  ram[39142]  = 1;
  ram[39143]  = 1;
  ram[39144]  = 1;
  ram[39145]  = 1;
  ram[39146]  = 1;
  ram[39147]  = 1;
  ram[39148]  = 1;
  ram[39149]  = 1;
  ram[39150]  = 1;
  ram[39151]  = 1;
  ram[39152]  = 1;
  ram[39153]  = 1;
  ram[39154]  = 1;
  ram[39155]  = 1;
  ram[39156]  = 1;
  ram[39157]  = 1;
  ram[39158]  = 1;
  ram[39159]  = 1;
  ram[39160]  = 1;
  ram[39161]  = 1;
  ram[39162]  = 1;
  ram[39163]  = 1;
  ram[39164]  = 1;
  ram[39165]  = 1;
  ram[39166]  = 1;
  ram[39167]  = 1;
  ram[39168]  = 1;
  ram[39169]  = 1;
  ram[39170]  = 1;
  ram[39171]  = 1;
  ram[39172]  = 1;
  ram[39173]  = 1;
  ram[39174]  = 1;
  ram[39175]  = 1;
  ram[39176]  = 1;
  ram[39177]  = 1;
  ram[39178]  = 1;
  ram[39179]  = 1;
  ram[39180]  = 1;
  ram[39181]  = 1;
  ram[39182]  = 1;
  ram[39183]  = 1;
  ram[39184]  = 1;
  ram[39185]  = 1;
  ram[39186]  = 1;
  ram[39187]  = 1;
  ram[39188]  = 1;
  ram[39189]  = 1;
  ram[39190]  = 1;
  ram[39191]  = 1;
  ram[39192]  = 1;
  ram[39193]  = 1;
  ram[39194]  = 1;
  ram[39195]  = 1;
  ram[39196]  = 1;
  ram[39197]  = 1;
  ram[39198]  = 1;
  ram[39199]  = 1;
  ram[39200]  = 1;
  ram[39201]  = 1;
  ram[39202]  = 1;
  ram[39203]  = 1;
  ram[39204]  = 1;
  ram[39205]  = 1;
  ram[39206]  = 1;
  ram[39207]  = 1;
  ram[39208]  = 1;
  ram[39209]  = 1;
  ram[39210]  = 1;
  ram[39211]  = 1;
  ram[39212]  = 1;
  ram[39213]  = 1;
  ram[39214]  = 1;
  ram[39215]  = 1;
  ram[39216]  = 1;
  ram[39217]  = 1;
  ram[39218]  = 1;
  ram[39219]  = 1;
  ram[39220]  = 1;
  ram[39221]  = 1;
  ram[39222]  = 1;
  ram[39223]  = 1;
  ram[39224]  = 1;
  ram[39225]  = 1;
  ram[39226]  = 1;
  ram[39227]  = 1;
  ram[39228]  = 1;
  ram[39229]  = 1;
  ram[39230]  = 1;
  ram[39231]  = 1;
  ram[39232]  = 1;
  ram[39233]  = 1;
  ram[39234]  = 1;
  ram[39235]  = 1;
  ram[39236]  = 1;
  ram[39237]  = 1;
  ram[39238]  = 1;
  ram[39239]  = 1;
  ram[39240]  = 1;
  ram[39241]  = 1;
  ram[39242]  = 1;
  ram[39243]  = 1;
  ram[39244]  = 1;
  ram[39245]  = 1;
  ram[39246]  = 1;
  ram[39247]  = 1;
  ram[39248]  = 1;
  ram[39249]  = 1;
  ram[39250]  = 1;
  ram[39251]  = 1;
  ram[39252]  = 1;
  ram[39253]  = 1;
  ram[39254]  = 1;
  ram[39255]  = 1;
  ram[39256]  = 1;
  ram[39257]  = 1;
  ram[39258]  = 1;
  ram[39259]  = 1;
  ram[39260]  = 1;
  ram[39261]  = 1;
  ram[39262]  = 1;
  ram[39263]  = 1;
  ram[39264]  = 1;
  ram[39265]  = 1;
  ram[39266]  = 1;
  ram[39267]  = 1;
  ram[39268]  = 1;
  ram[39269]  = 1;
  ram[39270]  = 1;
  ram[39271]  = 1;
  ram[39272]  = 1;
  ram[39273]  = 1;
  ram[39274]  = 1;
  ram[39275]  = 1;
  ram[39276]  = 1;
  ram[39277]  = 1;
  ram[39278]  = 1;
  ram[39279]  = 1;
  ram[39280]  = 1;
  ram[39281]  = 1;
  ram[39282]  = 1;
  ram[39283]  = 1;
  ram[39284]  = 1;
  ram[39285]  = 1;
  ram[39286]  = 1;
  ram[39287]  = 1;
  ram[39288]  = 1;
  ram[39289]  = 1;
  ram[39290]  = 1;
  ram[39291]  = 1;
  ram[39292]  = 1;
  ram[39293]  = 1;
  ram[39294]  = 1;
  ram[39295]  = 1;
  ram[39296]  = 1;
  ram[39297]  = 1;
  ram[39298]  = 1;
  ram[39299]  = 1;
  ram[39300]  = 1;
  ram[39301]  = 1;
  ram[39302]  = 1;
  ram[39303]  = 1;
  ram[39304]  = 1;
  ram[39305]  = 1;
  ram[39306]  = 1;
  ram[39307]  = 1;
  ram[39308]  = 1;
  ram[39309]  = 1;
  ram[39310]  = 1;
  ram[39311]  = 1;
  ram[39312]  = 1;
  ram[39313]  = 1;
  ram[39314]  = 1;
  ram[39315]  = 1;
  ram[39316]  = 1;
  ram[39317]  = 1;
  ram[39318]  = 1;
  ram[39319]  = 1;
  ram[39320]  = 1;
  ram[39321]  = 1;
  ram[39322]  = 1;
  ram[39323]  = 1;
  ram[39324]  = 1;
  ram[39325]  = 1;
  ram[39326]  = 1;
  ram[39327]  = 1;
  ram[39328]  = 1;
  ram[39329]  = 1;
  ram[39330]  = 1;
  ram[39331]  = 1;
  ram[39332]  = 1;
  ram[39333]  = 1;
  ram[39334]  = 1;
  ram[39335]  = 1;
  ram[39336]  = 1;
  ram[39337]  = 1;
  ram[39338]  = 1;
  ram[39339]  = 1;
  ram[39340]  = 1;
  ram[39341]  = 1;
  ram[39342]  = 1;
  ram[39343]  = 1;
  ram[39344]  = 1;
  ram[39345]  = 1;
  ram[39346]  = 1;
  ram[39347]  = 1;
  ram[39348]  = 1;
  ram[39349]  = 1;
  ram[39350]  = 1;
  ram[39351]  = 1;
  ram[39352]  = 1;
  ram[39353]  = 1;
  ram[39354]  = 1;
  ram[39355]  = 1;
  ram[39356]  = 1;
  ram[39357]  = 1;
  ram[39358]  = 1;
  ram[39359]  = 1;
  ram[39360]  = 1;
  ram[39361]  = 1;
  ram[39362]  = 1;
  ram[39363]  = 1;
  ram[39364]  = 1;
  ram[39365]  = 1;
  ram[39366]  = 1;
  ram[39367]  = 1;
  ram[39368]  = 1;
  ram[39369]  = 1;
  ram[39370]  = 1;
  ram[39371]  = 1;
  ram[39372]  = 1;
  ram[39373]  = 1;
  ram[39374]  = 1;
  ram[39375]  = 1;
  ram[39376]  = 1;
  ram[39377]  = 1;
  ram[39378]  = 1;
  ram[39379]  = 1;
  ram[39380]  = 1;
  ram[39381]  = 1;
  ram[39382]  = 1;
  ram[39383]  = 1;
  ram[39384]  = 1;
  ram[39385]  = 1;
  ram[39386]  = 1;
  ram[39387]  = 1;
  ram[39388]  = 1;
  ram[39389]  = 1;
  ram[39390]  = 1;
  ram[39391]  = 1;
  ram[39392]  = 1;
  ram[39393]  = 1;
  ram[39394]  = 1;
  ram[39395]  = 1;
  ram[39396]  = 1;
  ram[39397]  = 1;
  ram[39398]  = 1;
  ram[39399]  = 1;
  ram[39400]  = 1;
  ram[39401]  = 1;
  ram[39402]  = 1;
  ram[39403]  = 1;
  ram[39404]  = 1;
  ram[39405]  = 1;
  ram[39406]  = 1;
  ram[39407]  = 1;
  ram[39408]  = 1;
  ram[39409]  = 1;
  ram[39410]  = 1;
  ram[39411]  = 1;
  ram[39412]  = 1;
  ram[39413]  = 1;
  ram[39414]  = 1;
  ram[39415]  = 1;
  ram[39416]  = 1;
  ram[39417]  = 1;
  ram[39418]  = 1;
  ram[39419]  = 1;
  ram[39420]  = 1;
  ram[39421]  = 1;
  ram[39422]  = 1;
  ram[39423]  = 1;
  ram[39424]  = 1;
  ram[39425]  = 1;
  ram[39426]  = 1;
  ram[39427]  = 1;
  ram[39428]  = 1;
  ram[39429]  = 1;
  ram[39430]  = 1;
  ram[39431]  = 1;
  ram[39432]  = 1;
  ram[39433]  = 1;
  ram[39434]  = 1;
  ram[39435]  = 1;
  ram[39436]  = 1;
  ram[39437]  = 1;
  ram[39438]  = 1;
  ram[39439]  = 1;
  ram[39440]  = 1;
  ram[39441]  = 1;
  ram[39442]  = 1;
  ram[39443]  = 1;
  ram[39444]  = 1;
  ram[39445]  = 1;
  ram[39446]  = 1;
  ram[39447]  = 1;
  ram[39448]  = 1;
  ram[39449]  = 1;
  ram[39450]  = 1;
  ram[39451]  = 1;
  ram[39452]  = 1;
  ram[39453]  = 1;
  ram[39454]  = 1;
  ram[39455]  = 1;
  ram[39456]  = 1;
  ram[39457]  = 1;
  ram[39458]  = 1;
  ram[39459]  = 1;
  ram[39460]  = 1;
  ram[39461]  = 1;
  ram[39462]  = 1;
  ram[39463]  = 1;
  ram[39464]  = 1;
  ram[39465]  = 1;
  ram[39466]  = 1;
  ram[39467]  = 1;
  ram[39468]  = 1;
  ram[39469]  = 1;
  ram[39470]  = 1;
  ram[39471]  = 1;
  ram[39472]  = 1;
  ram[39473]  = 1;
  ram[39474]  = 1;
  ram[39475]  = 1;
  ram[39476]  = 1;
  ram[39477]  = 1;
  ram[39478]  = 1;
  ram[39479]  = 1;
  ram[39480]  = 1;
  ram[39481]  = 1;
  ram[39482]  = 1;
  ram[39483]  = 1;
  ram[39484]  = 1;
  ram[39485]  = 1;
  ram[39486]  = 1;
  ram[39487]  = 1;
  ram[39488]  = 1;
  ram[39489]  = 1;
  ram[39490]  = 1;
  ram[39491]  = 1;
  ram[39492]  = 1;
  ram[39493]  = 1;
  ram[39494]  = 1;
  ram[39495]  = 1;
  ram[39496]  = 1;
  ram[39497]  = 1;
  ram[39498]  = 1;
  ram[39499]  = 1;
  ram[39500]  = 1;
  ram[39501]  = 1;
  ram[39502]  = 1;
  ram[39503]  = 1;
  ram[39504]  = 1;
  ram[39505]  = 1;
  ram[39506]  = 1;
  ram[39507]  = 1;
  ram[39508]  = 1;
  ram[39509]  = 1;
  ram[39510]  = 1;
  ram[39511]  = 1;
  ram[39512]  = 1;
  ram[39513]  = 1;
  ram[39514]  = 1;
  ram[39515]  = 1;
  ram[39516]  = 1;
  ram[39517]  = 1;
  ram[39518]  = 1;
  ram[39519]  = 1;
  ram[39520]  = 1;
  ram[39521]  = 1;
  ram[39522]  = 1;
  ram[39523]  = 1;
  ram[39524]  = 1;
  ram[39525]  = 1;
  ram[39526]  = 1;
  ram[39527]  = 1;
  ram[39528]  = 1;
  ram[39529]  = 1;
  ram[39530]  = 1;
  ram[39531]  = 1;
  ram[39532]  = 1;
  ram[39533]  = 1;
  ram[39534]  = 1;
  ram[39535]  = 1;
  ram[39536]  = 1;
  ram[39537]  = 1;
  ram[39538]  = 1;
  ram[39539]  = 1;
  ram[39540]  = 1;
  ram[39541]  = 1;
  ram[39542]  = 1;
  ram[39543]  = 1;
  ram[39544]  = 1;
  ram[39545]  = 1;
  ram[39546]  = 1;
  ram[39547]  = 1;
  ram[39548]  = 1;
  ram[39549]  = 1;
  ram[39550]  = 1;
  ram[39551]  = 1;
  ram[39552]  = 1;
  ram[39553]  = 1;
  ram[39554]  = 1;
  ram[39555]  = 1;
  ram[39556]  = 1;
  ram[39557]  = 1;
  ram[39558]  = 1;
  ram[39559]  = 1;
  ram[39560]  = 1;
  ram[39561]  = 1;
  ram[39562]  = 1;
  ram[39563]  = 1;
  ram[39564]  = 1;
  ram[39565]  = 1;
  ram[39566]  = 1;
  ram[39567]  = 1;
  ram[39568]  = 1;
  ram[39569]  = 1;
  ram[39570]  = 1;
  ram[39571]  = 1;
  ram[39572]  = 1;
  ram[39573]  = 1;
  ram[39574]  = 1;
  ram[39575]  = 1;
  ram[39576]  = 1;
  ram[39577]  = 1;
  ram[39578]  = 1;
  ram[39579]  = 1;
  ram[39580]  = 1;
  ram[39581]  = 1;
  ram[39582]  = 1;
  ram[39583]  = 1;
  ram[39584]  = 1;
  ram[39585]  = 1;
  ram[39586]  = 1;
  ram[39587]  = 1;
  ram[39588]  = 1;
  ram[39589]  = 1;
  ram[39590]  = 1;
  ram[39591]  = 1;
  ram[39592]  = 1;
  ram[39593]  = 1;
  ram[39594]  = 1;
  ram[39595]  = 1;
  ram[39596]  = 1;
  ram[39597]  = 1;
  ram[39598]  = 1;
  ram[39599]  = 1;
  ram[39600]  = 1;
  ram[39601]  = 1;
  ram[39602]  = 1;
  ram[39603]  = 1;
  ram[39604]  = 1;
  ram[39605]  = 1;
  ram[39606]  = 1;
  ram[39607]  = 1;
  ram[39608]  = 1;
  ram[39609]  = 1;
  ram[39610]  = 1;
  ram[39611]  = 1;
  ram[39612]  = 1;
  ram[39613]  = 1;
  ram[39614]  = 1;
  ram[39615]  = 1;
  ram[39616]  = 1;
  ram[39617]  = 1;
  ram[39618]  = 1;
  ram[39619]  = 1;
  ram[39620]  = 1;
  ram[39621]  = 1;
  ram[39622]  = 1;
  ram[39623]  = 1;
  ram[39624]  = 1;
  ram[39625]  = 1;
  ram[39626]  = 1;
  ram[39627]  = 1;
  ram[39628]  = 1;
  ram[39629]  = 1;
  ram[39630]  = 1;
  ram[39631]  = 1;
  ram[39632]  = 1;
  ram[39633]  = 1;
  ram[39634]  = 1;
  ram[39635]  = 1;
  ram[39636]  = 1;
  ram[39637]  = 1;
  ram[39638]  = 1;
  ram[39639]  = 1;
  ram[39640]  = 1;
  ram[39641]  = 1;
  ram[39642]  = 1;
  ram[39643]  = 1;
  ram[39644]  = 1;
  ram[39645]  = 1;
  ram[39646]  = 1;
  ram[39647]  = 1;
  ram[39648]  = 1;
  ram[39649]  = 1;
  ram[39650]  = 1;
  ram[39651]  = 1;
  ram[39652]  = 1;
  ram[39653]  = 1;
  ram[39654]  = 1;
  ram[39655]  = 1;
  ram[39656]  = 1;
  ram[39657]  = 1;
  ram[39658]  = 1;
  ram[39659]  = 1;
  ram[39660]  = 1;
  ram[39661]  = 1;
  ram[39662]  = 1;
  ram[39663]  = 1;
  ram[39664]  = 1;
  ram[39665]  = 1;
  ram[39666]  = 1;
  ram[39667]  = 1;
  ram[39668]  = 1;
  ram[39669]  = 1;
  ram[39670]  = 1;
  ram[39671]  = 1;
  ram[39672]  = 1;
  ram[39673]  = 1;
  ram[39674]  = 1;
  ram[39675]  = 1;
  ram[39676]  = 1;
  ram[39677]  = 1;
  ram[39678]  = 1;
  ram[39679]  = 1;
  ram[39680]  = 1;
  ram[39681]  = 1;
  ram[39682]  = 1;
  ram[39683]  = 1;
  ram[39684]  = 1;
  ram[39685]  = 1;
  ram[39686]  = 1;
  ram[39687]  = 1;
  ram[39688]  = 1;
  ram[39689]  = 1;
  ram[39690]  = 1;
  ram[39691]  = 1;
  ram[39692]  = 1;
  ram[39693]  = 1;
  ram[39694]  = 1;
  ram[39695]  = 1;
  ram[39696]  = 1;
  ram[39697]  = 1;
  ram[39698]  = 1;
  ram[39699]  = 1;
  ram[39700]  = 1;
  ram[39701]  = 1;
  ram[39702]  = 1;
  ram[39703]  = 1;
  ram[39704]  = 1;
  ram[39705]  = 1;
  ram[39706]  = 1;
  ram[39707]  = 1;
  ram[39708]  = 1;
  ram[39709]  = 1;
  ram[39710]  = 1;
  ram[39711]  = 1;
  ram[39712]  = 1;
  ram[39713]  = 1;
  ram[39714]  = 1;
  ram[39715]  = 1;
  ram[39716]  = 1;
  ram[39717]  = 1;
  ram[39718]  = 1;
  ram[39719]  = 1;
  ram[39720]  = 1;
  ram[39721]  = 1;
  ram[39722]  = 1;
  ram[39723]  = 1;
  ram[39724]  = 1;
  ram[39725]  = 1;
  ram[39726]  = 1;
  ram[39727]  = 1;
  ram[39728]  = 1;
  ram[39729]  = 1;
  ram[39730]  = 1;
  ram[39731]  = 1;
  ram[39732]  = 1;
  ram[39733]  = 1;
  ram[39734]  = 1;
  ram[39735]  = 1;
  ram[39736]  = 1;
  ram[39737]  = 1;
  ram[39738]  = 1;
  ram[39739]  = 1;
  ram[39740]  = 1;
  ram[39741]  = 1;
  ram[39742]  = 1;
  ram[39743]  = 1;
  ram[39744]  = 1;
  ram[39745]  = 1;
  ram[39746]  = 1;
  ram[39747]  = 1;
  ram[39748]  = 1;
  ram[39749]  = 1;
  ram[39750]  = 1;
  ram[39751]  = 1;
  ram[39752]  = 1;
  ram[39753]  = 1;
  ram[39754]  = 1;
  ram[39755]  = 1;
  ram[39756]  = 1;
  ram[39757]  = 1;
  ram[39758]  = 1;
  ram[39759]  = 1;
  ram[39760]  = 1;
  ram[39761]  = 1;
  ram[39762]  = 1;
  ram[39763]  = 1;
  ram[39764]  = 1;
  ram[39765]  = 1;
  ram[39766]  = 1;
  ram[39767]  = 1;
  ram[39768]  = 1;
  ram[39769]  = 1;
  ram[39770]  = 1;
  ram[39771]  = 1;
  ram[39772]  = 1;
  ram[39773]  = 1;
  ram[39774]  = 1;
  ram[39775]  = 1;
  ram[39776]  = 1;
  ram[39777]  = 1;
  ram[39778]  = 1;
  ram[39779]  = 1;
  ram[39780]  = 1;
  ram[39781]  = 1;
  ram[39782]  = 1;
  ram[39783]  = 1;
  ram[39784]  = 1;
  ram[39785]  = 1;
  ram[39786]  = 1;
  ram[39787]  = 1;
  ram[39788]  = 1;
  ram[39789]  = 1;
  ram[39790]  = 1;
  ram[39791]  = 1;
  ram[39792]  = 1;
  ram[39793]  = 1;
  ram[39794]  = 1;
  ram[39795]  = 1;
  ram[39796]  = 1;
  ram[39797]  = 1;
  ram[39798]  = 1;
  ram[39799]  = 1;
  ram[39800]  = 1;
  ram[39801]  = 1;
  ram[39802]  = 1;
  ram[39803]  = 1;
  ram[39804]  = 1;
  ram[39805]  = 1;
  ram[39806]  = 1;
  ram[39807]  = 1;
  ram[39808]  = 1;
  ram[39809]  = 1;
  ram[39810]  = 1;
  ram[39811]  = 1;
  ram[39812]  = 1;
  ram[39813]  = 1;
  ram[39814]  = 1;
  ram[39815]  = 1;
  ram[39816]  = 1;
  ram[39817]  = 1;
  ram[39818]  = 1;
  ram[39819]  = 1;
  ram[39820]  = 1;
  ram[39821]  = 1;
  ram[39822]  = 1;
  ram[39823]  = 1;
  ram[39824]  = 1;
  ram[39825]  = 1;
  ram[39826]  = 1;
  ram[39827]  = 1;
  ram[39828]  = 1;
  ram[39829]  = 1;
  ram[39830]  = 1;
  ram[39831]  = 1;
  ram[39832]  = 1;
  ram[39833]  = 1;
  ram[39834]  = 1;
  ram[39835]  = 1;
  ram[39836]  = 1;
  ram[39837]  = 1;
  ram[39838]  = 1;
  ram[39839]  = 1;
  ram[39840]  = 1;
  ram[39841]  = 1;
  ram[39842]  = 1;
  ram[39843]  = 1;
  ram[39844]  = 1;
  ram[39845]  = 1;
  ram[39846]  = 1;
  ram[39847]  = 1;
  ram[39848]  = 1;
  ram[39849]  = 1;
  ram[39850]  = 1;
  ram[39851]  = 1;
  ram[39852]  = 1;
  ram[39853]  = 1;
  ram[39854]  = 1;
  ram[39855]  = 1;
  ram[39856]  = 1;
  ram[39857]  = 1;
  ram[39858]  = 1;
  ram[39859]  = 1;
  ram[39860]  = 1;
  ram[39861]  = 1;
  ram[39862]  = 1;
  ram[39863]  = 1;
  ram[39864]  = 1;
  ram[39865]  = 1;
  ram[39866]  = 1;
  ram[39867]  = 1;
  ram[39868]  = 1;
  ram[39869]  = 1;
  ram[39870]  = 1;
  ram[39871]  = 1;
  ram[39872]  = 1;
  ram[39873]  = 1;
  ram[39874]  = 1;
  ram[39875]  = 1;
  ram[39876]  = 1;
  ram[39877]  = 1;
  ram[39878]  = 1;
  ram[39879]  = 1;
  ram[39880]  = 1;
  ram[39881]  = 1;
  ram[39882]  = 1;
  ram[39883]  = 1;
  ram[39884]  = 1;
  ram[39885]  = 1;
  ram[39886]  = 1;
  ram[39887]  = 1;
  ram[39888]  = 1;
  ram[39889]  = 1;
  ram[39890]  = 1;
  ram[39891]  = 1;
  ram[39892]  = 1;
  ram[39893]  = 1;
  ram[39894]  = 1;
  ram[39895]  = 1;
  ram[39896]  = 1;
  ram[39897]  = 1;
  ram[39898]  = 1;
  ram[39899]  = 1;
  ram[39900]  = 1;
  ram[39901]  = 1;
  ram[39902]  = 1;
  ram[39903]  = 1;
  ram[39904]  = 1;
  ram[39905]  = 1;
  ram[39906]  = 1;
  ram[39907]  = 1;
  ram[39908]  = 1;
  ram[39909]  = 1;
  ram[39910]  = 1;
  ram[39911]  = 1;
  ram[39912]  = 1;
  ram[39913]  = 1;
  ram[39914]  = 1;
  ram[39915]  = 1;
  ram[39916]  = 1;
  ram[39917]  = 1;
  ram[39918]  = 1;
  ram[39919]  = 1;
  ram[39920]  = 1;
  ram[39921]  = 1;
  ram[39922]  = 1;
  ram[39923]  = 1;
  ram[39924]  = 1;
  ram[39925]  = 1;
  ram[39926]  = 1;
  ram[39927]  = 1;
  ram[39928]  = 1;
  ram[39929]  = 1;
  ram[39930]  = 1;
  ram[39931]  = 1;
  ram[39932]  = 1;
  ram[39933]  = 1;
  ram[39934]  = 1;
  ram[39935]  = 1;
  ram[39936]  = 1;
  ram[39937]  = 1;
  ram[39938]  = 1;
  ram[39939]  = 1;
  ram[39940]  = 1;
  ram[39941]  = 1;
  ram[39942]  = 1;
  ram[39943]  = 1;
  ram[39944]  = 1;
  ram[39945]  = 1;
  ram[39946]  = 1;
  ram[39947]  = 1;
  ram[39948]  = 1;
  ram[39949]  = 1;
  ram[39950]  = 1;
  ram[39951]  = 1;
  ram[39952]  = 1;
  ram[39953]  = 1;
  ram[39954]  = 1;
  ram[39955]  = 1;
  ram[39956]  = 1;
  ram[39957]  = 1;
  ram[39958]  = 1;
  ram[39959]  = 1;
  ram[39960]  = 1;
  ram[39961]  = 1;
  ram[39962]  = 1;
  ram[39963]  = 1;
  ram[39964]  = 1;
  ram[39965]  = 1;
  ram[39966]  = 1;
  ram[39967]  = 1;
  ram[39968]  = 1;
  ram[39969]  = 1;
  ram[39970]  = 1;
  ram[39971]  = 1;
  ram[39972]  = 1;
  ram[39973]  = 1;
  ram[39974]  = 1;
  ram[39975]  = 1;
  ram[39976]  = 1;
  ram[39977]  = 1;
  ram[39978]  = 1;
  ram[39979]  = 1;
  ram[39980]  = 1;
  ram[39981]  = 1;
  ram[39982]  = 1;
  ram[39983]  = 1;
  ram[39984]  = 1;
  ram[39985]  = 1;
  ram[39986]  = 1;
  ram[39987]  = 1;
  ram[39988]  = 1;
  ram[39989]  = 1;
  ram[39990]  = 1;
  ram[39991]  = 1;
  ram[39992]  = 1;
  ram[39993]  = 1;
  ram[39994]  = 1;
  ram[39995]  = 1;
  ram[39996]  = 1;
  ram[39997]  = 1;
  ram[39998]  = 1;
  ram[39999]  = 1;
  ram[40000]  = 1;
  ram[40001]  = 1;
  ram[40002]  = 1;
  ram[40003]  = 1;
  ram[40004]  = 1;
  ram[40005]  = 1;
  ram[40006]  = 1;
  ram[40007]  = 1;
  ram[40008]  = 1;
  ram[40009]  = 1;
  ram[40010]  = 1;
  ram[40011]  = 1;
  ram[40012]  = 1;
  ram[40013]  = 1;
  ram[40014]  = 1;
  ram[40015]  = 1;
  ram[40016]  = 1;
  ram[40017]  = 1;
  ram[40018]  = 1;
  ram[40019]  = 1;
  ram[40020]  = 1;
  ram[40021]  = 1;
  ram[40022]  = 1;
  ram[40023]  = 1;
  ram[40024]  = 1;
  ram[40025]  = 1;
  ram[40026]  = 1;
  ram[40027]  = 1;
  ram[40028]  = 1;
  ram[40029]  = 1;
  ram[40030]  = 1;
  ram[40031]  = 1;
  ram[40032]  = 1;
  ram[40033]  = 1;
  ram[40034]  = 1;
  ram[40035]  = 1;
  ram[40036]  = 1;
  ram[40037]  = 1;
  ram[40038]  = 1;
  ram[40039]  = 1;
  ram[40040]  = 1;
  ram[40041]  = 1;
  ram[40042]  = 1;
  ram[40043]  = 1;
  ram[40044]  = 1;
  ram[40045]  = 1;
  ram[40046]  = 1;
  ram[40047]  = 1;
  ram[40048]  = 1;
  ram[40049]  = 1;
  ram[40050]  = 1;
  ram[40051]  = 1;
  ram[40052]  = 1;
  ram[40053]  = 1;
  ram[40054]  = 1;
  ram[40055]  = 1;
  ram[40056]  = 1;
  ram[40057]  = 1;
  ram[40058]  = 1;
  ram[40059]  = 1;
  ram[40060]  = 1;
  ram[40061]  = 1;
  ram[40062]  = 1;
  ram[40063]  = 1;
  ram[40064]  = 1;
  ram[40065]  = 1;
  ram[40066]  = 1;
  ram[40067]  = 1;
  ram[40068]  = 1;
  ram[40069]  = 1;
  ram[40070]  = 1;
  ram[40071]  = 1;
  ram[40072]  = 1;
  ram[40073]  = 1;
  ram[40074]  = 1;
  ram[40075]  = 1;
  ram[40076]  = 1;
  ram[40077]  = 1;
  ram[40078]  = 1;
  ram[40079]  = 1;
  ram[40080]  = 1;
  ram[40081]  = 1;
  ram[40082]  = 1;
  ram[40083]  = 1;
  ram[40084]  = 1;
  ram[40085]  = 1;
  ram[40086]  = 1;
  ram[40087]  = 1;
  ram[40088]  = 1;
  ram[40089]  = 1;
  ram[40090]  = 1;
  ram[40091]  = 1;
  ram[40092]  = 1;
  ram[40093]  = 1;
  ram[40094]  = 1;
  ram[40095]  = 1;
  ram[40096]  = 1;
  ram[40097]  = 1;
  ram[40098]  = 1;
  ram[40099]  = 1;
  ram[40100]  = 1;
  ram[40101]  = 1;
  ram[40102]  = 1;
  ram[40103]  = 1;
  ram[40104]  = 1;
  ram[40105]  = 1;
  ram[40106]  = 1;
  ram[40107]  = 1;
  ram[40108]  = 1;
  ram[40109]  = 1;
  ram[40110]  = 1;
  ram[40111]  = 1;
  ram[40112]  = 1;
  ram[40113]  = 1;
  ram[40114]  = 1;
  ram[40115]  = 1;
  ram[40116]  = 1;
  ram[40117]  = 1;
  ram[40118]  = 1;
  ram[40119]  = 1;
  ram[40120]  = 1;
  ram[40121]  = 1;
  ram[40122]  = 1;
  ram[40123]  = 1;
  ram[40124]  = 1;
  ram[40125]  = 1;
  ram[40126]  = 1;
  ram[40127]  = 1;
  ram[40128]  = 1;
  ram[40129]  = 1;
  ram[40130]  = 1;
  ram[40131]  = 1;
  ram[40132]  = 1;
  ram[40133]  = 1;
  ram[40134]  = 1;
  ram[40135]  = 1;
  ram[40136]  = 1;
  ram[40137]  = 1;
  ram[40138]  = 1;
  ram[40139]  = 1;
  ram[40140]  = 1;
  ram[40141]  = 1;
  ram[40142]  = 1;
  ram[40143]  = 1;
  ram[40144]  = 1;
  ram[40145]  = 1;
  ram[40146]  = 1;
  ram[40147]  = 1;
  ram[40148]  = 1;
  ram[40149]  = 1;
  ram[40150]  = 1;
  ram[40151]  = 1;
  ram[40152]  = 1;
  ram[40153]  = 1;
  ram[40154]  = 1;
  ram[40155]  = 1;
  ram[40156]  = 1;
  ram[40157]  = 1;
  ram[40158]  = 1;
  ram[40159]  = 1;
  ram[40160]  = 1;
  ram[40161]  = 1;
  ram[40162]  = 1;
  ram[40163]  = 1;
  ram[40164]  = 1;
  ram[40165]  = 1;
  ram[40166]  = 1;
  ram[40167]  = 1;
  ram[40168]  = 1;
  ram[40169]  = 1;
  ram[40170]  = 1;
  ram[40171]  = 1;
  ram[40172]  = 1;
  ram[40173]  = 1;
  ram[40174]  = 1;
  ram[40175]  = 1;
  ram[40176]  = 1;
  ram[40177]  = 1;
  ram[40178]  = 1;
  ram[40179]  = 1;
  ram[40180]  = 1;
  ram[40181]  = 1;
  ram[40182]  = 1;
  ram[40183]  = 1;
  ram[40184]  = 1;
  ram[40185]  = 1;
  ram[40186]  = 1;
  ram[40187]  = 1;
  ram[40188]  = 1;
  ram[40189]  = 1;
  ram[40190]  = 1;
  ram[40191]  = 1;
  ram[40192]  = 1;
  ram[40193]  = 1;
  ram[40194]  = 1;
  ram[40195]  = 1;
  ram[40196]  = 1;
  ram[40197]  = 1;
  ram[40198]  = 1;
  ram[40199]  = 1;
  ram[40200]  = 1;
  ram[40201]  = 1;
  ram[40202]  = 1;
  ram[40203]  = 1;
  ram[40204]  = 1;
  ram[40205]  = 1;
  ram[40206]  = 1;
  ram[40207]  = 1;
  ram[40208]  = 1;
  ram[40209]  = 1;
  ram[40210]  = 1;
  ram[40211]  = 1;
  ram[40212]  = 1;
  ram[40213]  = 1;
  ram[40214]  = 1;
  ram[40215]  = 1;
  ram[40216]  = 1;
  ram[40217]  = 1;
  ram[40218]  = 1;
  ram[40219]  = 1;
  ram[40220]  = 1;
  ram[40221]  = 1;
  ram[40222]  = 1;
  ram[40223]  = 1;
  ram[40224]  = 1;
  ram[40225]  = 1;
  ram[40226]  = 1;
  ram[40227]  = 1;
  ram[40228]  = 1;
  ram[40229]  = 1;
  ram[40230]  = 1;
  ram[40231]  = 1;
  ram[40232]  = 1;
  ram[40233]  = 1;
  ram[40234]  = 1;
  ram[40235]  = 1;
  ram[40236]  = 1;
  ram[40237]  = 1;
  ram[40238]  = 1;
  ram[40239]  = 1;
  ram[40240]  = 1;
  ram[40241]  = 1;
  ram[40242]  = 1;
  ram[40243]  = 1;
  ram[40244]  = 1;
  ram[40245]  = 1;
  ram[40246]  = 1;
  ram[40247]  = 1;
  ram[40248]  = 1;
  ram[40249]  = 1;
  ram[40250]  = 1;
  ram[40251]  = 1;
  ram[40252]  = 1;
  ram[40253]  = 1;
  ram[40254]  = 1;
  ram[40255]  = 1;
  ram[40256]  = 1;
  ram[40257]  = 1;
  ram[40258]  = 1;
  ram[40259]  = 1;
  ram[40260]  = 1;
  ram[40261]  = 1;
  ram[40262]  = 1;
  ram[40263]  = 1;
  ram[40264]  = 1;
  ram[40265]  = 1;
  ram[40266]  = 1;
  ram[40267]  = 1;
  ram[40268]  = 1;
  ram[40269]  = 1;
  ram[40270]  = 1;
  ram[40271]  = 1;
  ram[40272]  = 1;
  ram[40273]  = 1;
  ram[40274]  = 1;
  ram[40275]  = 1;
  ram[40276]  = 1;
  ram[40277]  = 1;
  ram[40278]  = 1;
  ram[40279]  = 1;
  ram[40280]  = 1;
  ram[40281]  = 1;
  ram[40282]  = 1;
  ram[40283]  = 1;
  ram[40284]  = 1;
  ram[40285]  = 1;
  ram[40286]  = 1;
  ram[40287]  = 1;
  ram[40288]  = 1;
  ram[40289]  = 1;
  ram[40290]  = 1;
  ram[40291]  = 1;
  ram[40292]  = 1;
  ram[40293]  = 1;
  ram[40294]  = 1;
  ram[40295]  = 1;
  ram[40296]  = 1;
  ram[40297]  = 1;
  ram[40298]  = 1;
  ram[40299]  = 1;
  ram[40300]  = 1;
  ram[40301]  = 1;
  ram[40302]  = 1;
  ram[40303]  = 1;
  ram[40304]  = 1;
  ram[40305]  = 1;
  ram[40306]  = 1;
  ram[40307]  = 1;
  ram[40308]  = 1;
  ram[40309]  = 1;
  ram[40310]  = 1;
  ram[40311]  = 1;
  ram[40312]  = 1;
  ram[40313]  = 1;
  ram[40314]  = 1;
  ram[40315]  = 1;
  ram[40316]  = 1;
  ram[40317]  = 1;
  ram[40318]  = 1;
  ram[40319]  = 1;
  ram[40320]  = 1;
  ram[40321]  = 1;
  ram[40322]  = 1;
  ram[40323]  = 1;
  ram[40324]  = 1;
  ram[40325]  = 1;
  ram[40326]  = 1;
  ram[40327]  = 1;
  ram[40328]  = 1;
  ram[40329]  = 1;
  ram[40330]  = 1;
  ram[40331]  = 1;
  ram[40332]  = 1;
  ram[40333]  = 1;
  ram[40334]  = 1;
  ram[40335]  = 1;
  ram[40336]  = 1;
  ram[40337]  = 1;
  ram[40338]  = 1;
  ram[40339]  = 1;
  ram[40340]  = 1;
  ram[40341]  = 1;
  ram[40342]  = 1;
  ram[40343]  = 1;
  ram[40344]  = 1;
  ram[40345]  = 1;
  ram[40346]  = 1;
  ram[40347]  = 1;
  ram[40348]  = 1;
  ram[40349]  = 1;
  ram[40350]  = 1;
  ram[40351]  = 1;
  ram[40352]  = 1;
  ram[40353]  = 1;
  ram[40354]  = 1;
  ram[40355]  = 1;
  ram[40356]  = 1;
  ram[40357]  = 1;
  ram[40358]  = 1;
  ram[40359]  = 1;
  ram[40360]  = 1;
  ram[40361]  = 1;
  ram[40362]  = 1;
  ram[40363]  = 1;
  ram[40364]  = 1;
  ram[40365]  = 1;
  ram[40366]  = 1;
  ram[40367]  = 1;
  ram[40368]  = 1;
  ram[40369]  = 1;
  ram[40370]  = 1;
  ram[40371]  = 1;
  ram[40372]  = 1;
  ram[40373]  = 1;
  ram[40374]  = 1;
  ram[40375]  = 1;
  ram[40376]  = 1;
  ram[40377]  = 1;
  ram[40378]  = 1;
  ram[40379]  = 1;
  ram[40380]  = 1;
  ram[40381]  = 1;
  ram[40382]  = 1;
  ram[40383]  = 1;
  ram[40384]  = 1;
  ram[40385]  = 1;
  ram[40386]  = 1;
  ram[40387]  = 1;
  ram[40388]  = 1;
  ram[40389]  = 1;
  ram[40390]  = 1;
  ram[40391]  = 1;
  ram[40392]  = 1;
  ram[40393]  = 1;
  ram[40394]  = 1;
  ram[40395]  = 1;
  ram[40396]  = 1;
  ram[40397]  = 1;
  ram[40398]  = 1;
  ram[40399]  = 1;
  ram[40400]  = 1;
  ram[40401]  = 1;
  ram[40402]  = 1;
  ram[40403]  = 1;
  ram[40404]  = 1;
  ram[40405]  = 1;
  ram[40406]  = 1;
  ram[40407]  = 1;
  ram[40408]  = 1;
  ram[40409]  = 1;
  ram[40410]  = 1;
  ram[40411]  = 1;
  ram[40412]  = 1;
  ram[40413]  = 1;
  ram[40414]  = 1;
  ram[40415]  = 1;
  ram[40416]  = 1;
  ram[40417]  = 1;
  ram[40418]  = 1;
  ram[40419]  = 1;
  ram[40420]  = 1;
  ram[40421]  = 1;
  ram[40422]  = 1;
  ram[40423]  = 1;
  ram[40424]  = 1;
  ram[40425]  = 1;
  ram[40426]  = 1;
  ram[40427]  = 1;
  ram[40428]  = 1;
  ram[40429]  = 1;
  ram[40430]  = 1;
  ram[40431]  = 1;
  ram[40432]  = 1;
  ram[40433]  = 1;
  ram[40434]  = 1;
  ram[40435]  = 1;
  ram[40436]  = 1;
  ram[40437]  = 1;
  ram[40438]  = 1;
  ram[40439]  = 1;
  ram[40440]  = 1;
  ram[40441]  = 1;
  ram[40442]  = 1;
  ram[40443]  = 1;
  ram[40444]  = 1;
  ram[40445]  = 1;
  ram[40446]  = 1;
  ram[40447]  = 1;
  ram[40448]  = 1;
  ram[40449]  = 1;
  ram[40450]  = 1;
  ram[40451]  = 1;
  ram[40452]  = 1;
  ram[40453]  = 1;
  ram[40454]  = 1;
  ram[40455]  = 1;
  ram[40456]  = 1;
  ram[40457]  = 1;
  ram[40458]  = 1;
  ram[40459]  = 1;
  ram[40460]  = 1;
  ram[40461]  = 1;
  ram[40462]  = 1;
  ram[40463]  = 1;
  ram[40464]  = 1;
  ram[40465]  = 1;
  ram[40466]  = 1;
  ram[40467]  = 1;
  ram[40468]  = 1;
  ram[40469]  = 1;
  ram[40470]  = 1;
  ram[40471]  = 1;
  ram[40472]  = 1;
  ram[40473]  = 1;
  ram[40474]  = 1;
  ram[40475]  = 1;
  ram[40476]  = 1;
  ram[40477]  = 1;
  ram[40478]  = 1;
  ram[40479]  = 1;
  ram[40480]  = 1;
  ram[40481]  = 1;
  ram[40482]  = 1;
  ram[40483]  = 1;
  ram[40484]  = 1;
  ram[40485]  = 1;
  ram[40486]  = 1;
  ram[40487]  = 1;
  ram[40488]  = 1;
  ram[40489]  = 1;
  ram[40490]  = 1;
  ram[40491]  = 1;
  ram[40492]  = 1;
  ram[40493]  = 1;
  ram[40494]  = 1;
  ram[40495]  = 1;
  ram[40496]  = 1;
  ram[40497]  = 1;
  ram[40498]  = 1;
  ram[40499]  = 1;
  ram[40500]  = 1;
  ram[40501]  = 1;
  ram[40502]  = 1;
  ram[40503]  = 1;
  ram[40504]  = 1;
  ram[40505]  = 1;
  ram[40506]  = 1;
  ram[40507]  = 1;
  ram[40508]  = 1;
  ram[40509]  = 1;
  ram[40510]  = 1;
  ram[40511]  = 1;
  ram[40512]  = 1;
  ram[40513]  = 1;
  ram[40514]  = 1;
  ram[40515]  = 1;
  ram[40516]  = 1;
  ram[40517]  = 1;
  ram[40518]  = 1;
  ram[40519]  = 1;
  ram[40520]  = 1;
  ram[40521]  = 1;
  ram[40522]  = 1;
  ram[40523]  = 1;
  ram[40524]  = 1;
  ram[40525]  = 1;
  ram[40526]  = 1;
  ram[40527]  = 1;
  ram[40528]  = 1;
  ram[40529]  = 1;
  ram[40530]  = 1;
  ram[40531]  = 1;
  ram[40532]  = 1;
  ram[40533]  = 1;
  ram[40534]  = 1;
  ram[40535]  = 1;
  ram[40536]  = 1;
  ram[40537]  = 1;
  ram[40538]  = 1;
  ram[40539]  = 1;
  ram[40540]  = 1;
  ram[40541]  = 1;
  ram[40542]  = 1;
  ram[40543]  = 1;
  ram[40544]  = 1;
  ram[40545]  = 1;
  ram[40546]  = 1;
  ram[40547]  = 1;
  ram[40548]  = 1;
  ram[40549]  = 1;
  ram[40550]  = 1;
  ram[40551]  = 1;
  ram[40552]  = 1;
  ram[40553]  = 1;
  ram[40554]  = 1;
  ram[40555]  = 1;
  ram[40556]  = 1;
  ram[40557]  = 1;
  ram[40558]  = 1;
  ram[40559]  = 1;
  ram[40560]  = 1;
  ram[40561]  = 1;
  ram[40562]  = 1;
  ram[40563]  = 1;
  ram[40564]  = 1;
  ram[40565]  = 1;
  ram[40566]  = 1;
  ram[40567]  = 1;
  ram[40568]  = 1;
  ram[40569]  = 1;
  ram[40570]  = 1;
  ram[40571]  = 1;
  ram[40572]  = 1;
  ram[40573]  = 1;
  ram[40574]  = 1;
  ram[40575]  = 1;
  ram[40576]  = 1;
  ram[40577]  = 1;
  ram[40578]  = 1;
  ram[40579]  = 1;
  ram[40580]  = 1;
  ram[40581]  = 1;
  ram[40582]  = 1;
  ram[40583]  = 1;
  ram[40584]  = 1;
  ram[40585]  = 1;
  ram[40586]  = 1;
  ram[40587]  = 1;
  ram[40588]  = 1;
  ram[40589]  = 1;
  ram[40590]  = 1;
  ram[40591]  = 1;
  ram[40592]  = 1;
  ram[40593]  = 1;
  ram[40594]  = 1;
  ram[40595]  = 1;
  ram[40596]  = 1;
  ram[40597]  = 1;
  ram[40598]  = 1;
  ram[40599]  = 1;
  ram[40600]  = 1;
  ram[40601]  = 1;
  ram[40602]  = 1;
  ram[40603]  = 1;
  ram[40604]  = 1;
  ram[40605]  = 1;
  ram[40606]  = 1;
  ram[40607]  = 1;
  ram[40608]  = 1;
  ram[40609]  = 1;
  ram[40610]  = 1;
  ram[40611]  = 1;
  ram[40612]  = 1;
  ram[40613]  = 1;
  ram[40614]  = 1;
  ram[40615]  = 1;
  ram[40616]  = 1;
  ram[40617]  = 1;
  ram[40618]  = 1;
  ram[40619]  = 1;
  ram[40620]  = 1;
  ram[40621]  = 1;
  ram[40622]  = 1;
  ram[40623]  = 1;
  ram[40624]  = 1;
  ram[40625]  = 1;
  ram[40626]  = 1;
  ram[40627]  = 1;
  ram[40628]  = 1;
  ram[40629]  = 1;
  ram[40630]  = 1;
  ram[40631]  = 1;
  ram[40632]  = 1;
  ram[40633]  = 1;
  ram[40634]  = 1;
  ram[40635]  = 1;
  ram[40636]  = 1;
  ram[40637]  = 1;
  ram[40638]  = 1;
  ram[40639]  = 1;
  ram[40640]  = 1;
  ram[40641]  = 1;
  ram[40642]  = 1;
  ram[40643]  = 1;
  ram[40644]  = 1;
  ram[40645]  = 1;
  ram[40646]  = 1;
  ram[40647]  = 1;
  ram[40648]  = 1;
  ram[40649]  = 1;
  ram[40650]  = 1;
  ram[40651]  = 1;
  ram[40652]  = 1;
  ram[40653]  = 1;
  ram[40654]  = 1;
  ram[40655]  = 1;
  ram[40656]  = 1;
  ram[40657]  = 1;
  ram[40658]  = 1;
  ram[40659]  = 1;
  ram[40660]  = 1;
  ram[40661]  = 1;
  ram[40662]  = 1;
  ram[40663]  = 1;
  ram[40664]  = 1;
  ram[40665]  = 1;
  ram[40666]  = 1;
  ram[40667]  = 1;
  ram[40668]  = 1;
  ram[40669]  = 1;
  ram[40670]  = 1;
  ram[40671]  = 1;
  ram[40672]  = 1;
  ram[40673]  = 1;
  ram[40674]  = 1;
  ram[40675]  = 1;
  ram[40676]  = 1;
  ram[40677]  = 1;
  ram[40678]  = 1;
  ram[40679]  = 1;
  ram[40680]  = 1;
  ram[40681]  = 1;
  ram[40682]  = 1;
  ram[40683]  = 1;
  ram[40684]  = 1;
  ram[40685]  = 1;
  ram[40686]  = 1;
  ram[40687]  = 1;
  ram[40688]  = 1;
  ram[40689]  = 1;
  ram[40690]  = 1;
  ram[40691]  = 1;
  ram[40692]  = 1;
  ram[40693]  = 1;
  ram[40694]  = 1;
  ram[40695]  = 1;
  ram[40696]  = 1;
  ram[40697]  = 1;
  ram[40698]  = 1;
  ram[40699]  = 1;
  ram[40700]  = 1;
  ram[40701]  = 1;
  ram[40702]  = 1;
  ram[40703]  = 1;
  ram[40704]  = 1;
  ram[40705]  = 1;
  ram[40706]  = 1;
  ram[40707]  = 1;
  ram[40708]  = 1;
  ram[40709]  = 1;
  ram[40710]  = 1;
  ram[40711]  = 1;
  ram[40712]  = 1;
  ram[40713]  = 1;
  ram[40714]  = 1;
  ram[40715]  = 1;
  ram[40716]  = 1;
  ram[40717]  = 1;
  ram[40718]  = 1;
  ram[40719]  = 1;
  ram[40720]  = 1;
  ram[40721]  = 1;
  ram[40722]  = 1;
  ram[40723]  = 1;
  ram[40724]  = 1;
  ram[40725]  = 1;
  ram[40726]  = 1;
  ram[40727]  = 1;
  ram[40728]  = 1;
  ram[40729]  = 1;
  ram[40730]  = 1;
  ram[40731]  = 1;
  ram[40732]  = 1;
  ram[40733]  = 1;
  ram[40734]  = 1;
  ram[40735]  = 1;
  ram[40736]  = 1;
  ram[40737]  = 1;
  ram[40738]  = 1;
  ram[40739]  = 1;
  ram[40740]  = 1;
  ram[40741]  = 1;
  ram[40742]  = 1;
  ram[40743]  = 1;
  ram[40744]  = 1;
  ram[40745]  = 1;
  ram[40746]  = 1;
  ram[40747]  = 1;
  ram[40748]  = 1;
  ram[40749]  = 1;
  ram[40750]  = 1;
  ram[40751]  = 1;
  ram[40752]  = 1;
  ram[40753]  = 1;
  ram[40754]  = 1;
  ram[40755]  = 1;
  ram[40756]  = 1;
  ram[40757]  = 1;
  ram[40758]  = 1;
  ram[40759]  = 1;
  ram[40760]  = 1;
  ram[40761]  = 1;
  ram[40762]  = 1;
  ram[40763]  = 1;
  ram[40764]  = 1;
  ram[40765]  = 1;
  ram[40766]  = 1;
  ram[40767]  = 1;
  ram[40768]  = 1;
  ram[40769]  = 1;
  ram[40770]  = 1;
  ram[40771]  = 1;
  ram[40772]  = 1;
  ram[40773]  = 1;
  ram[40774]  = 1;
  ram[40775]  = 1;
  ram[40776]  = 1;
  ram[40777]  = 1;
  ram[40778]  = 1;
  ram[40779]  = 1;
  ram[40780]  = 1;
  ram[40781]  = 1;
  ram[40782]  = 1;
  ram[40783]  = 1;
  ram[40784]  = 1;
  ram[40785]  = 1;
  ram[40786]  = 1;
  ram[40787]  = 1;
  ram[40788]  = 1;
  ram[40789]  = 1;
  ram[40790]  = 1;
  ram[40791]  = 1;
  ram[40792]  = 1;
  ram[40793]  = 1;
  ram[40794]  = 1;
  ram[40795]  = 1;
  ram[40796]  = 1;
  ram[40797]  = 1;
  ram[40798]  = 1;
  ram[40799]  = 1;
  ram[40800]  = 1;
  ram[40801]  = 1;
  ram[40802]  = 1;
  ram[40803]  = 1;
  ram[40804]  = 1;
  ram[40805]  = 1;
  ram[40806]  = 1;
  ram[40807]  = 1;
  ram[40808]  = 1;
  ram[40809]  = 1;
  ram[40810]  = 1;
  ram[40811]  = 1;
  ram[40812]  = 1;
  ram[40813]  = 1;
  ram[40814]  = 1;
  ram[40815]  = 1;
  ram[40816]  = 1;
  ram[40817]  = 1;
  ram[40818]  = 1;
  ram[40819]  = 1;
  ram[40820]  = 1;
  ram[40821]  = 1;
  ram[40822]  = 1;
  ram[40823]  = 1;
  ram[40824]  = 1;
  ram[40825]  = 1;
  ram[40826]  = 1;
  ram[40827]  = 1;
  ram[40828]  = 1;
  ram[40829]  = 1;
  ram[40830]  = 1;
  ram[40831]  = 1;
  ram[40832]  = 1;
  ram[40833]  = 1;
  ram[40834]  = 1;
  ram[40835]  = 1;
  ram[40836]  = 1;
  ram[40837]  = 1;
  ram[40838]  = 1;
  ram[40839]  = 1;
  ram[40840]  = 1;
  ram[40841]  = 1;
  ram[40842]  = 1;
  ram[40843]  = 1;
  ram[40844]  = 1;
  ram[40845]  = 1;
  ram[40846]  = 1;
  ram[40847]  = 1;
  ram[40848]  = 1;
  ram[40849]  = 1;
  ram[40850]  = 1;
  ram[40851]  = 1;
  ram[40852]  = 1;
  ram[40853]  = 1;
  ram[40854]  = 1;
  ram[40855]  = 1;
  ram[40856]  = 1;
  ram[40857]  = 1;
  ram[40858]  = 1;
  ram[40859]  = 1;
  ram[40860]  = 1;
  ram[40861]  = 1;
  ram[40862]  = 1;
  ram[40863]  = 1;
  ram[40864]  = 1;
  ram[40865]  = 1;
  ram[40866]  = 1;
  ram[40867]  = 1;
  ram[40868]  = 1;
  ram[40869]  = 1;
  ram[40870]  = 1;
  ram[40871]  = 1;
  ram[40872]  = 1;
  ram[40873]  = 1;
  ram[40874]  = 1;
  ram[40875]  = 1;
  ram[40876]  = 1;
  ram[40877]  = 1;
  ram[40878]  = 1;
  ram[40879]  = 1;
  ram[40880]  = 1;
  ram[40881]  = 1;
  ram[40882]  = 1;
  ram[40883]  = 1;
  ram[40884]  = 1;
  ram[40885]  = 1;
  ram[40886]  = 1;
  ram[40887]  = 1;
  ram[40888]  = 1;
  ram[40889]  = 1;
  ram[40890]  = 1;
  ram[40891]  = 1;
  ram[40892]  = 1;
  ram[40893]  = 1;
  ram[40894]  = 1;
  ram[40895]  = 1;
  ram[40896]  = 1;
  ram[40897]  = 1;
  ram[40898]  = 1;
  ram[40899]  = 1;
  ram[40900]  = 1;
  ram[40901]  = 1;
  ram[40902]  = 1;
  ram[40903]  = 1;
  ram[40904]  = 1;
  ram[40905]  = 1;
  ram[40906]  = 1;
  ram[40907]  = 1;
  ram[40908]  = 1;
  ram[40909]  = 1;
  ram[40910]  = 1;
  ram[40911]  = 1;
  ram[40912]  = 1;
  ram[40913]  = 1;
  ram[40914]  = 1;
  ram[40915]  = 1;
  ram[40916]  = 1;
  ram[40917]  = 1;
  ram[40918]  = 1;
  ram[40919]  = 1;
  ram[40920]  = 1;
  ram[40921]  = 1;
  ram[40922]  = 1;
  ram[40923]  = 1;
  ram[40924]  = 1;
  ram[40925]  = 1;
  ram[40926]  = 1;
  ram[40927]  = 1;
  ram[40928]  = 1;
  ram[40929]  = 1;
  ram[40930]  = 1;
  ram[40931]  = 1;
  ram[40932]  = 1;
  ram[40933]  = 1;
  ram[40934]  = 1;
  ram[40935]  = 1;
  ram[40936]  = 1;
  ram[40937]  = 1;
  ram[40938]  = 1;
  ram[40939]  = 1;
  ram[40940]  = 1;
  ram[40941]  = 1;
  ram[40942]  = 1;
  ram[40943]  = 1;
  ram[40944]  = 1;
  ram[40945]  = 1;
  ram[40946]  = 1;
  ram[40947]  = 1;
  ram[40948]  = 1;
  ram[40949]  = 1;
  ram[40950]  = 1;
  ram[40951]  = 1;
  ram[40952]  = 1;
  ram[40953]  = 1;
  ram[40954]  = 1;
  ram[40955]  = 1;
  ram[40956]  = 1;
  ram[40957]  = 1;
  ram[40958]  = 1;
  ram[40959]  = 1;
  ram[40960]  = 1;
  ram[40961]  = 1;
  ram[40962]  = 1;
  ram[40963]  = 1;
  ram[40964]  = 1;
  ram[40965]  = 1;
  ram[40966]  = 1;
  ram[40967]  = 1;
  ram[40968]  = 1;
  ram[40969]  = 1;
  ram[40970]  = 1;
  ram[40971]  = 1;
  ram[40972]  = 1;
  ram[40973]  = 1;
  ram[40974]  = 1;
  ram[40975]  = 1;
  ram[40976]  = 1;
  ram[40977]  = 1;
  ram[40978]  = 1;
  ram[40979]  = 1;
  ram[40980]  = 1;
  ram[40981]  = 1;
  ram[40982]  = 1;
  ram[40983]  = 1;
  ram[40984]  = 1;
  ram[40985]  = 1;
  ram[40986]  = 1;
  ram[40987]  = 1;
  ram[40988]  = 1;
  ram[40989]  = 1;
  ram[40990]  = 1;
  ram[40991]  = 1;
  ram[40992]  = 1;
  ram[40993]  = 1;
  ram[40994]  = 1;
  ram[40995]  = 1;
  ram[40996]  = 1;
  ram[40997]  = 1;
  ram[40998]  = 1;
  ram[40999]  = 1;
  ram[41000]  = 1;
  ram[41001]  = 1;
  ram[41002]  = 1;
  ram[41003]  = 1;
  ram[41004]  = 1;
  ram[41005]  = 1;
  ram[41006]  = 1;
  ram[41007]  = 1;
  ram[41008]  = 1;
  ram[41009]  = 1;
  ram[41010]  = 1;
  ram[41011]  = 1;
  ram[41012]  = 1;
  ram[41013]  = 1;
  ram[41014]  = 1;
  ram[41015]  = 1;
  ram[41016]  = 1;
  ram[41017]  = 1;
  ram[41018]  = 1;
  ram[41019]  = 1;
  ram[41020]  = 1;
  ram[41021]  = 1;
  ram[41022]  = 1;
  ram[41023]  = 1;
  ram[41024]  = 1;
  ram[41025]  = 1;
  ram[41026]  = 1;
  ram[41027]  = 1;
  ram[41028]  = 1;
  ram[41029]  = 1;
  ram[41030]  = 1;
  ram[41031]  = 1;
  ram[41032]  = 1;
  ram[41033]  = 1;
  ram[41034]  = 1;
  ram[41035]  = 1;
  ram[41036]  = 1;
  ram[41037]  = 1;
  ram[41038]  = 1;
  ram[41039]  = 1;
  ram[41040]  = 1;
  ram[41041]  = 1;
  ram[41042]  = 1;
  ram[41043]  = 1;
  ram[41044]  = 1;
  ram[41045]  = 1;
  ram[41046]  = 1;
  ram[41047]  = 1;
  ram[41048]  = 1;
  ram[41049]  = 1;
  ram[41050]  = 1;
  ram[41051]  = 1;
  ram[41052]  = 1;
  ram[41053]  = 1;
  ram[41054]  = 1;
  ram[41055]  = 1;
  ram[41056]  = 1;
  ram[41057]  = 1;
  ram[41058]  = 1;
  ram[41059]  = 1;
  ram[41060]  = 1;
  ram[41061]  = 1;
  ram[41062]  = 1;
  ram[41063]  = 1;
  ram[41064]  = 1;
  ram[41065]  = 1;
  ram[41066]  = 1;
  ram[41067]  = 1;
  ram[41068]  = 1;
  ram[41069]  = 1;
  ram[41070]  = 1;
  ram[41071]  = 1;
  ram[41072]  = 1;
  ram[41073]  = 1;
  ram[41074]  = 1;
  ram[41075]  = 1;
  ram[41076]  = 1;
  ram[41077]  = 1;
  ram[41078]  = 1;
  ram[41079]  = 1;
  ram[41080]  = 1;
  ram[41081]  = 1;
  ram[41082]  = 1;
  ram[41083]  = 1;
  ram[41084]  = 1;
  ram[41085]  = 1;
  ram[41086]  = 1;
  ram[41087]  = 1;
  ram[41088]  = 1;
  ram[41089]  = 1;
  ram[41090]  = 1;
  ram[41091]  = 1;
  ram[41092]  = 1;
  ram[41093]  = 1;
  ram[41094]  = 1;
  ram[41095]  = 1;
  ram[41096]  = 1;
  ram[41097]  = 1;
  ram[41098]  = 1;
  ram[41099]  = 1;
  ram[41100]  = 1;
  ram[41101]  = 1;
  ram[41102]  = 1;
  ram[41103]  = 1;
  ram[41104]  = 1;
  ram[41105]  = 1;
  ram[41106]  = 1;
  ram[41107]  = 1;
  ram[41108]  = 1;
  ram[41109]  = 1;
  ram[41110]  = 1;
  ram[41111]  = 1;
  ram[41112]  = 1;
  ram[41113]  = 1;
  ram[41114]  = 1;
  ram[41115]  = 1;
  ram[41116]  = 1;
  ram[41117]  = 1;
  ram[41118]  = 1;
  ram[41119]  = 1;
  ram[41120]  = 1;
  ram[41121]  = 1;
  ram[41122]  = 1;
  ram[41123]  = 1;
  ram[41124]  = 1;
  ram[41125]  = 1;
  ram[41126]  = 1;
  ram[41127]  = 1;
  ram[41128]  = 1;
  ram[41129]  = 1;
  ram[41130]  = 1;
  ram[41131]  = 1;
  ram[41132]  = 1;
  ram[41133]  = 1;
  ram[41134]  = 1;
  ram[41135]  = 1;
  ram[41136]  = 1;
  ram[41137]  = 1;
  ram[41138]  = 1;
  ram[41139]  = 1;
  ram[41140]  = 1;
  ram[41141]  = 1;
  ram[41142]  = 1;
  ram[41143]  = 1;
  ram[41144]  = 1;
  ram[41145]  = 1;
  ram[41146]  = 1;
  ram[41147]  = 1;
  ram[41148]  = 1;
  ram[41149]  = 1;
  ram[41150]  = 1;
  ram[41151]  = 1;
  ram[41152]  = 1;
  ram[41153]  = 1;
  ram[41154]  = 1;
  ram[41155]  = 1;
  ram[41156]  = 1;
  ram[41157]  = 1;
  ram[41158]  = 1;
  ram[41159]  = 1;
  ram[41160]  = 1;
  ram[41161]  = 1;
  ram[41162]  = 1;
  ram[41163]  = 1;
  ram[41164]  = 1;
  ram[41165]  = 1;
  ram[41166]  = 1;
  ram[41167]  = 1;
  ram[41168]  = 1;
  ram[41169]  = 1;
  ram[41170]  = 1;
  ram[41171]  = 1;
  ram[41172]  = 1;
  ram[41173]  = 1;
  ram[41174]  = 1;
  ram[41175]  = 1;
  ram[41176]  = 1;
  ram[41177]  = 1;
  ram[41178]  = 1;
  ram[41179]  = 1;
  ram[41180]  = 1;
  ram[41181]  = 1;
  ram[41182]  = 1;
  ram[41183]  = 1;
  ram[41184]  = 1;
  ram[41185]  = 1;
  ram[41186]  = 1;
  ram[41187]  = 1;
  ram[41188]  = 1;
  ram[41189]  = 1;
  ram[41190]  = 1;
  ram[41191]  = 1;
  ram[41192]  = 1;
  ram[41193]  = 1;
  ram[41194]  = 1;
  ram[41195]  = 1;
  ram[41196]  = 1;
  ram[41197]  = 1;
  ram[41198]  = 1;
  ram[41199]  = 1;
  ram[41200]  = 1;
  ram[41201]  = 1;
  ram[41202]  = 1;
  ram[41203]  = 1;
  ram[41204]  = 1;
  ram[41205]  = 1;
  ram[41206]  = 1;
  ram[41207]  = 1;
  ram[41208]  = 1;
  ram[41209]  = 1;
  ram[41210]  = 1;
  ram[41211]  = 1;
  ram[41212]  = 1;
  ram[41213]  = 1;
  ram[41214]  = 1;
  ram[41215]  = 1;
  ram[41216]  = 1;
  ram[41217]  = 1;
  ram[41218]  = 1;
  ram[41219]  = 1;
  ram[41220]  = 1;
  ram[41221]  = 1;
  ram[41222]  = 1;
  ram[41223]  = 1;
  ram[41224]  = 1;
  ram[41225]  = 1;
  ram[41226]  = 1;
  ram[41227]  = 1;
  ram[41228]  = 1;
  ram[41229]  = 1;
  ram[41230]  = 1;
  ram[41231]  = 1;
  ram[41232]  = 1;
  ram[41233]  = 1;
  ram[41234]  = 1;
  ram[41235]  = 1;
  ram[41236]  = 1;
  ram[41237]  = 1;
  ram[41238]  = 1;
  ram[41239]  = 1;
  ram[41240]  = 1;
  ram[41241]  = 1;
  ram[41242]  = 1;
  ram[41243]  = 1;
  ram[41244]  = 1;
  ram[41245]  = 1;
  ram[41246]  = 1;
  ram[41247]  = 1;
  ram[41248]  = 1;
  ram[41249]  = 1;
  ram[41250]  = 1;
  ram[41251]  = 1;
  ram[41252]  = 1;
  ram[41253]  = 1;
  ram[41254]  = 1;
  ram[41255]  = 1;
  ram[41256]  = 1;
  ram[41257]  = 1;
  ram[41258]  = 1;
  ram[41259]  = 1;
  ram[41260]  = 1;
  ram[41261]  = 1;
  ram[41262]  = 1;
  ram[41263]  = 1;
  ram[41264]  = 1;
  ram[41265]  = 1;
  ram[41266]  = 1;
  ram[41267]  = 1;
  ram[41268]  = 1;
  ram[41269]  = 1;
  ram[41270]  = 1;
  ram[41271]  = 1;
  ram[41272]  = 1;
  ram[41273]  = 1;
  ram[41274]  = 1;
  ram[41275]  = 1;
  ram[41276]  = 1;
  ram[41277]  = 1;
  ram[41278]  = 1;
  ram[41279]  = 1;
  ram[41280]  = 1;
  ram[41281]  = 1;
  ram[41282]  = 1;
  ram[41283]  = 1;
  ram[41284]  = 1;
  ram[41285]  = 1;
  ram[41286]  = 1;
  ram[41287]  = 1;
  ram[41288]  = 1;
  ram[41289]  = 1;
  ram[41290]  = 1;
  ram[41291]  = 1;
  ram[41292]  = 1;
  ram[41293]  = 1;
  ram[41294]  = 1;
  ram[41295]  = 1;
  ram[41296]  = 1;
  ram[41297]  = 1;
  ram[41298]  = 1;
  ram[41299]  = 1;
  ram[41300]  = 1;
  ram[41301]  = 1;
  ram[41302]  = 1;
  ram[41303]  = 1;
  ram[41304]  = 1;
  ram[41305]  = 1;
  ram[41306]  = 1;
  ram[41307]  = 1;
  ram[41308]  = 1;
  ram[41309]  = 1;
  ram[41310]  = 1;
  ram[41311]  = 1;
  ram[41312]  = 1;
  ram[41313]  = 1;
  ram[41314]  = 1;
  ram[41315]  = 1;
  ram[41316]  = 1;
  ram[41317]  = 1;
  ram[41318]  = 1;
  ram[41319]  = 1;
  ram[41320]  = 1;
  ram[41321]  = 1;
  ram[41322]  = 1;
  ram[41323]  = 1;
  ram[41324]  = 1;
  ram[41325]  = 1;
  ram[41326]  = 1;
  ram[41327]  = 1;
  ram[41328]  = 1;
  ram[41329]  = 1;
  ram[41330]  = 1;
  ram[41331]  = 1;
  ram[41332]  = 1;
  ram[41333]  = 1;
  ram[41334]  = 1;
  ram[41335]  = 1;
  ram[41336]  = 1;
  ram[41337]  = 1;
  ram[41338]  = 1;
  ram[41339]  = 1;
  ram[41340]  = 1;
  ram[41341]  = 1;
  ram[41342]  = 1;
  ram[41343]  = 1;
  ram[41344]  = 1;
  ram[41345]  = 1;
  ram[41346]  = 1;
  ram[41347]  = 1;
  ram[41348]  = 1;
  ram[41349]  = 1;
  ram[41350]  = 1;
  ram[41351]  = 1;
  ram[41352]  = 1;
  ram[41353]  = 1;
  ram[41354]  = 1;
  ram[41355]  = 1;
  ram[41356]  = 1;
  ram[41357]  = 1;
  ram[41358]  = 1;
  ram[41359]  = 1;
  ram[41360]  = 1;
  ram[41361]  = 1;
  ram[41362]  = 1;
  ram[41363]  = 1;
  ram[41364]  = 1;
  ram[41365]  = 1;
  ram[41366]  = 1;
  ram[41367]  = 1;
  ram[41368]  = 1;
  ram[41369]  = 1;
  ram[41370]  = 1;
  ram[41371]  = 1;
  ram[41372]  = 1;
  ram[41373]  = 1;
  ram[41374]  = 1;
  ram[41375]  = 1;
  ram[41376]  = 1;
  ram[41377]  = 1;
  ram[41378]  = 1;
  ram[41379]  = 1;
  ram[41380]  = 1;
  ram[41381]  = 1;
  ram[41382]  = 1;
  ram[41383]  = 1;
  ram[41384]  = 1;
  ram[41385]  = 1;
  ram[41386]  = 1;
  ram[41387]  = 1;
  ram[41388]  = 1;
  ram[41389]  = 1;
  ram[41390]  = 1;
  ram[41391]  = 1;
  ram[41392]  = 1;
  ram[41393]  = 1;
  ram[41394]  = 1;
  ram[41395]  = 1;
  ram[41396]  = 1;
  ram[41397]  = 1;
  ram[41398]  = 1;
  ram[41399]  = 1;
  ram[41400]  = 1;
  ram[41401]  = 1;
  ram[41402]  = 1;
  ram[41403]  = 1;
  ram[41404]  = 1;
  ram[41405]  = 1;
  ram[41406]  = 1;
  ram[41407]  = 1;
  ram[41408]  = 1;
  ram[41409]  = 1;
  ram[41410]  = 1;
  ram[41411]  = 1;
  ram[41412]  = 1;
  ram[41413]  = 1;
  ram[41414]  = 1;
  ram[41415]  = 1;
  ram[41416]  = 1;
  ram[41417]  = 1;
  ram[41418]  = 1;
  ram[41419]  = 1;
  ram[41420]  = 1;
  ram[41421]  = 1;
  ram[41422]  = 1;
  ram[41423]  = 1;
  ram[41424]  = 1;
  ram[41425]  = 1;
  ram[41426]  = 1;
  ram[41427]  = 1;
  ram[41428]  = 1;
  ram[41429]  = 1;
  ram[41430]  = 1;
  ram[41431]  = 1;
  ram[41432]  = 1;
  ram[41433]  = 1;
  ram[41434]  = 1;
  ram[41435]  = 1;
  ram[41436]  = 1;
  ram[41437]  = 1;
  ram[41438]  = 1;
  ram[41439]  = 1;
  ram[41440]  = 1;
  ram[41441]  = 1;
  ram[41442]  = 1;
  ram[41443]  = 1;
  ram[41444]  = 1;
  ram[41445]  = 1;
  ram[41446]  = 1;
  ram[41447]  = 1;
  ram[41448]  = 1;
  ram[41449]  = 1;
  ram[41450]  = 1;
  ram[41451]  = 1;
  ram[41452]  = 1;
  ram[41453]  = 1;
  ram[41454]  = 1;
  ram[41455]  = 1;
  ram[41456]  = 1;
  ram[41457]  = 1;
  ram[41458]  = 1;
  ram[41459]  = 1;
  ram[41460]  = 1;
  ram[41461]  = 1;
  ram[41462]  = 1;
  ram[41463]  = 1;
  ram[41464]  = 1;
  ram[41465]  = 1;
  ram[41466]  = 1;
  ram[41467]  = 1;
  ram[41468]  = 1;
  ram[41469]  = 1;
  ram[41470]  = 1;
  ram[41471]  = 1;
  ram[41472]  = 1;
  ram[41473]  = 1;
  ram[41474]  = 1;
  ram[41475]  = 1;
  ram[41476]  = 1;
  ram[41477]  = 1;
  ram[41478]  = 1;
  ram[41479]  = 1;
  ram[41480]  = 1;
  ram[41481]  = 1;
  ram[41482]  = 1;
  ram[41483]  = 1;
  ram[41484]  = 1;
  ram[41485]  = 1;
  ram[41486]  = 1;
  ram[41487]  = 1;
  ram[41488]  = 1;
  ram[41489]  = 1;
  ram[41490]  = 1;
  ram[41491]  = 1;
  ram[41492]  = 1;
  ram[41493]  = 1;
  ram[41494]  = 1;
  ram[41495]  = 1;
  ram[41496]  = 1;
  ram[41497]  = 1;
  ram[41498]  = 1;
  ram[41499]  = 1;
  ram[41500]  = 1;
  ram[41501]  = 1;
  ram[41502]  = 1;
  ram[41503]  = 1;
  ram[41504]  = 1;
  ram[41505]  = 1;
  ram[41506]  = 1;
  ram[41507]  = 1;
  ram[41508]  = 1;
  ram[41509]  = 1;
  ram[41510]  = 1;
  ram[41511]  = 1;
  ram[41512]  = 1;
  ram[41513]  = 1;
  ram[41514]  = 1;
  ram[41515]  = 1;
  ram[41516]  = 1;
  ram[41517]  = 1;
  ram[41518]  = 1;
  ram[41519]  = 1;
  ram[41520]  = 1;
  ram[41521]  = 1;
  ram[41522]  = 1;
  ram[41523]  = 1;
  ram[41524]  = 1;
  ram[41525]  = 1;
  ram[41526]  = 1;
  ram[41527]  = 1;
  ram[41528]  = 1;
  ram[41529]  = 1;
  ram[41530]  = 1;
  ram[41531]  = 1;
  ram[41532]  = 1;
  ram[41533]  = 1;
  ram[41534]  = 1;
  ram[41535]  = 1;
  ram[41536]  = 1;
  ram[41537]  = 1;
  ram[41538]  = 1;
  ram[41539]  = 1;
  ram[41540]  = 1;
  ram[41541]  = 1;
  ram[41542]  = 1;
  ram[41543]  = 1;
  ram[41544]  = 1;
  ram[41545]  = 1;
  ram[41546]  = 1;
  ram[41547]  = 1;
  ram[41548]  = 1;
  ram[41549]  = 1;
  ram[41550]  = 1;
  ram[41551]  = 1;
  ram[41552]  = 1;
  ram[41553]  = 1;
  ram[41554]  = 1;
  ram[41555]  = 1;
  ram[41556]  = 1;
  ram[41557]  = 1;
  ram[41558]  = 1;
  ram[41559]  = 1;
  ram[41560]  = 1;
  ram[41561]  = 1;
  ram[41562]  = 1;
  ram[41563]  = 1;
  ram[41564]  = 1;
  ram[41565]  = 1;
  ram[41566]  = 1;
  ram[41567]  = 1;
  ram[41568]  = 1;
  ram[41569]  = 1;
  ram[41570]  = 1;
  ram[41571]  = 1;
  ram[41572]  = 1;
  ram[41573]  = 1;
  ram[41574]  = 1;
  ram[41575]  = 1;
  ram[41576]  = 1;
  ram[41577]  = 1;
  ram[41578]  = 1;
  ram[41579]  = 1;
  ram[41580]  = 1;
  ram[41581]  = 1;
  ram[41582]  = 1;
  ram[41583]  = 1;
  ram[41584]  = 1;
  ram[41585]  = 1;
  ram[41586]  = 1;
  ram[41587]  = 1;
  ram[41588]  = 1;
  ram[41589]  = 1;
  ram[41590]  = 1;
  ram[41591]  = 1;
  ram[41592]  = 1;
  ram[41593]  = 1;
  ram[41594]  = 1;
  ram[41595]  = 1;
  ram[41596]  = 1;
  ram[41597]  = 1;
  ram[41598]  = 1;
  ram[41599]  = 1;
  ram[41600]  = 1;
  ram[41601]  = 1;
  ram[41602]  = 1;
  ram[41603]  = 1;
  ram[41604]  = 1;
  ram[41605]  = 1;
  ram[41606]  = 1;
  ram[41607]  = 1;
  ram[41608]  = 1;
  ram[41609]  = 1;
  ram[41610]  = 1;
  ram[41611]  = 1;
  ram[41612]  = 1;
  ram[41613]  = 1;
  ram[41614]  = 1;
  ram[41615]  = 1;
  ram[41616]  = 1;
  ram[41617]  = 1;
  ram[41618]  = 1;
  ram[41619]  = 1;
  ram[41620]  = 1;
  ram[41621]  = 1;
  ram[41622]  = 1;
  ram[41623]  = 1;
  ram[41624]  = 1;
  ram[41625]  = 1;
  ram[41626]  = 1;
  ram[41627]  = 1;
  ram[41628]  = 1;
  ram[41629]  = 1;
  ram[41630]  = 1;
  ram[41631]  = 1;
  ram[41632]  = 1;
  ram[41633]  = 1;
  ram[41634]  = 1;
  ram[41635]  = 1;
  ram[41636]  = 1;
  ram[41637]  = 1;
  ram[41638]  = 1;
  ram[41639]  = 1;
  ram[41640]  = 1;
  ram[41641]  = 1;
  ram[41642]  = 1;
  ram[41643]  = 1;
  ram[41644]  = 1;
  ram[41645]  = 1;
  ram[41646]  = 1;
  ram[41647]  = 1;
  ram[41648]  = 1;
  ram[41649]  = 1;
  ram[41650]  = 1;
  ram[41651]  = 1;
  ram[41652]  = 1;
  ram[41653]  = 1;
  ram[41654]  = 1;
  ram[41655]  = 1;
  ram[41656]  = 1;
  ram[41657]  = 1;
  ram[41658]  = 1;
  ram[41659]  = 1;
  ram[41660]  = 1;
  ram[41661]  = 1;
  ram[41662]  = 1;
  ram[41663]  = 1;
  ram[41664]  = 1;
  ram[41665]  = 1;
  ram[41666]  = 1;
  ram[41667]  = 1;
  ram[41668]  = 1;
  ram[41669]  = 1;
  ram[41670]  = 1;
  ram[41671]  = 1;
  ram[41672]  = 1;
  ram[41673]  = 1;
  ram[41674]  = 1;
  ram[41675]  = 1;
  ram[41676]  = 1;
  ram[41677]  = 1;
  ram[41678]  = 1;
  ram[41679]  = 1;
  ram[41680]  = 1;
  ram[41681]  = 1;
  ram[41682]  = 1;
  ram[41683]  = 1;
  ram[41684]  = 1;
  ram[41685]  = 1;
  ram[41686]  = 1;
  ram[41687]  = 1;
  ram[41688]  = 1;
  ram[41689]  = 1;
  ram[41690]  = 1;
  ram[41691]  = 1;
  ram[41692]  = 1;
  ram[41693]  = 1;
  ram[41694]  = 1;
  ram[41695]  = 1;
  ram[41696]  = 1;
  ram[41697]  = 1;
  ram[41698]  = 1;
  ram[41699]  = 1;
  ram[41700]  = 1;
  ram[41701]  = 1;
  ram[41702]  = 1;
  ram[41703]  = 1;
  ram[41704]  = 1;
  ram[41705]  = 1;
  ram[41706]  = 1;
  ram[41707]  = 1;
  ram[41708]  = 1;
  ram[41709]  = 1;
  ram[41710]  = 1;
  ram[41711]  = 1;
  ram[41712]  = 1;
  ram[41713]  = 1;
  ram[41714]  = 1;
  ram[41715]  = 1;
  ram[41716]  = 1;
  ram[41717]  = 1;
  ram[41718]  = 1;
  ram[41719]  = 1;
  ram[41720]  = 1;
  ram[41721]  = 1;
  ram[41722]  = 1;
  ram[41723]  = 1;
  ram[41724]  = 1;
  ram[41725]  = 1;
  ram[41726]  = 1;
  ram[41727]  = 1;
  ram[41728]  = 1;
  ram[41729]  = 1;
  ram[41730]  = 1;
  ram[41731]  = 1;
  ram[41732]  = 1;
  ram[41733]  = 1;
  ram[41734]  = 1;
  ram[41735]  = 1;
  ram[41736]  = 1;
  ram[41737]  = 1;
  ram[41738]  = 1;
  ram[41739]  = 1;
  ram[41740]  = 1;
  ram[41741]  = 1;
  ram[41742]  = 1;
  ram[41743]  = 1;
  ram[41744]  = 1;
  ram[41745]  = 1;
  ram[41746]  = 1;
  ram[41747]  = 1;
  ram[41748]  = 1;
  ram[41749]  = 1;
  ram[41750]  = 1;
  ram[41751]  = 1;
  ram[41752]  = 1;
  ram[41753]  = 1;
  ram[41754]  = 1;
  ram[41755]  = 1;
  ram[41756]  = 1;
  ram[41757]  = 1;
  ram[41758]  = 1;
  ram[41759]  = 1;
  ram[41760]  = 1;
  ram[41761]  = 1;
  ram[41762]  = 1;
  ram[41763]  = 1;
  ram[41764]  = 1;
  ram[41765]  = 1;
  ram[41766]  = 1;
  ram[41767]  = 1;
  ram[41768]  = 1;
  ram[41769]  = 1;
  ram[41770]  = 1;
  ram[41771]  = 1;
  ram[41772]  = 1;
  ram[41773]  = 1;
  ram[41774]  = 1;
  ram[41775]  = 1;
  ram[41776]  = 1;
  ram[41777]  = 1;
  ram[41778]  = 1;
  ram[41779]  = 1;
  ram[41780]  = 1;
  ram[41781]  = 1;
  ram[41782]  = 1;
  ram[41783]  = 1;
  ram[41784]  = 1;
  ram[41785]  = 1;
  ram[41786]  = 1;
  ram[41787]  = 1;
  ram[41788]  = 1;
  ram[41789]  = 1;
  ram[41790]  = 1;
  ram[41791]  = 1;
  ram[41792]  = 1;
  ram[41793]  = 1;
  ram[41794]  = 1;
  ram[41795]  = 1;
  ram[41796]  = 1;
  ram[41797]  = 1;
  ram[41798]  = 1;
  ram[41799]  = 1;
  ram[41800]  = 1;
  ram[41801]  = 1;
  ram[41802]  = 1;
  ram[41803]  = 1;
  ram[41804]  = 1;
  ram[41805]  = 1;
  ram[41806]  = 1;
  ram[41807]  = 1;
  ram[41808]  = 1;
  ram[41809]  = 1;
  ram[41810]  = 1;
  ram[41811]  = 1;
  ram[41812]  = 1;
  ram[41813]  = 1;
  ram[41814]  = 1;
  ram[41815]  = 1;
  ram[41816]  = 1;
  ram[41817]  = 1;
  ram[41818]  = 1;
  ram[41819]  = 1;
  ram[41820]  = 1;
  ram[41821]  = 1;
  ram[41822]  = 1;
  ram[41823]  = 1;
  ram[41824]  = 1;
  ram[41825]  = 1;
  ram[41826]  = 1;
  ram[41827]  = 1;
  ram[41828]  = 1;
  ram[41829]  = 1;
  ram[41830]  = 1;
  ram[41831]  = 1;
  ram[41832]  = 1;
  ram[41833]  = 1;
  ram[41834]  = 1;
  ram[41835]  = 1;
  ram[41836]  = 1;
  ram[41837]  = 1;
  ram[41838]  = 1;
  ram[41839]  = 1;
  ram[41840]  = 1;
  ram[41841]  = 1;
  ram[41842]  = 1;
  ram[41843]  = 1;
  ram[41844]  = 1;
  ram[41845]  = 1;
  ram[41846]  = 1;
  ram[41847]  = 1;
  ram[41848]  = 1;
  ram[41849]  = 1;
  ram[41850]  = 1;
  ram[41851]  = 1;
  ram[41852]  = 1;
  ram[41853]  = 1;
  ram[41854]  = 1;
  ram[41855]  = 1;
  ram[41856]  = 1;
  ram[41857]  = 1;
  ram[41858]  = 1;
  ram[41859]  = 1;
  ram[41860]  = 1;
  ram[41861]  = 1;
  ram[41862]  = 1;
  ram[41863]  = 1;
  ram[41864]  = 1;
  ram[41865]  = 1;
  ram[41866]  = 1;
  ram[41867]  = 1;
  ram[41868]  = 1;
  ram[41869]  = 1;
  ram[41870]  = 1;
  ram[41871]  = 1;
  ram[41872]  = 1;
  ram[41873]  = 1;
  ram[41874]  = 1;
  ram[41875]  = 1;
  ram[41876]  = 1;
  ram[41877]  = 1;
  ram[41878]  = 1;
  ram[41879]  = 1;
  ram[41880]  = 1;
  ram[41881]  = 1;
  ram[41882]  = 1;
  ram[41883]  = 1;
  ram[41884]  = 1;
  ram[41885]  = 1;
  ram[41886]  = 1;
  ram[41887]  = 1;
  ram[41888]  = 1;
  ram[41889]  = 1;
  ram[41890]  = 1;
  ram[41891]  = 1;
  ram[41892]  = 1;
  ram[41893]  = 1;
  ram[41894]  = 1;
  ram[41895]  = 1;
  ram[41896]  = 1;
  ram[41897]  = 1;
  ram[41898]  = 1;
  ram[41899]  = 1;
  ram[41900]  = 1;
  ram[41901]  = 1;
  ram[41902]  = 1;
  ram[41903]  = 1;
  ram[41904]  = 1;
  ram[41905]  = 1;
  ram[41906]  = 1;
  ram[41907]  = 1;
  ram[41908]  = 1;
  ram[41909]  = 1;
  ram[41910]  = 1;
  ram[41911]  = 1;
  ram[41912]  = 1;
  ram[41913]  = 1;
  ram[41914]  = 1;
  ram[41915]  = 1;
  ram[41916]  = 1;
  ram[41917]  = 1;
  ram[41918]  = 1;
  ram[41919]  = 1;
  ram[41920]  = 1;
  ram[41921]  = 1;
  ram[41922]  = 1;
  ram[41923]  = 1;
  ram[41924]  = 1;
  ram[41925]  = 1;
  ram[41926]  = 1;
  ram[41927]  = 1;
  ram[41928]  = 1;
  ram[41929]  = 1;
  ram[41930]  = 1;
  ram[41931]  = 1;
  ram[41932]  = 1;
  ram[41933]  = 1;
  ram[41934]  = 1;
  ram[41935]  = 1;
  ram[41936]  = 1;
  ram[41937]  = 1;
  ram[41938]  = 1;
  ram[41939]  = 1;
  ram[41940]  = 1;
  ram[41941]  = 1;
  ram[41942]  = 1;
  ram[41943]  = 1;
  ram[41944]  = 1;
  ram[41945]  = 1;
  ram[41946]  = 1;
  ram[41947]  = 1;
  ram[41948]  = 1;
  ram[41949]  = 1;
  ram[41950]  = 1;
  ram[41951]  = 1;
  ram[41952]  = 1;
  ram[41953]  = 1;
  ram[41954]  = 1;
  ram[41955]  = 1;
  ram[41956]  = 1;
  ram[41957]  = 1;
  ram[41958]  = 1;
  ram[41959]  = 1;
  ram[41960]  = 1;
  ram[41961]  = 1;
  ram[41962]  = 1;
  ram[41963]  = 1;
  ram[41964]  = 1;
  ram[41965]  = 1;
  ram[41966]  = 1;
  ram[41967]  = 1;
  ram[41968]  = 1;
  ram[41969]  = 1;
  ram[41970]  = 1;
  ram[41971]  = 1;
  ram[41972]  = 1;
  ram[41973]  = 1;
  ram[41974]  = 1;
  ram[41975]  = 1;
  ram[41976]  = 1;
  ram[41977]  = 1;
  ram[41978]  = 1;
  ram[41979]  = 1;
  ram[41980]  = 1;
  ram[41981]  = 1;
  ram[41982]  = 1;
  ram[41983]  = 1;
  ram[41984]  = 1;
  ram[41985]  = 1;
  ram[41986]  = 1;
  ram[41987]  = 1;
  ram[41988]  = 1;
  ram[41989]  = 1;
  ram[41990]  = 1;
  ram[41991]  = 1;
  ram[41992]  = 1;
  ram[41993]  = 1;
  ram[41994]  = 1;
  ram[41995]  = 1;
  ram[41996]  = 1;
  ram[41997]  = 1;
  ram[41998]  = 1;
  ram[41999]  = 1;
  ram[42000]  = 1;
  ram[42001]  = 1;
  ram[42002]  = 1;
  ram[42003]  = 1;
  ram[42004]  = 1;
  ram[42005]  = 1;
  ram[42006]  = 1;
  ram[42007]  = 1;
  ram[42008]  = 1;
  ram[42009]  = 1;
  ram[42010]  = 1;
  ram[42011]  = 1;
  ram[42012]  = 1;
  ram[42013]  = 1;
  ram[42014]  = 1;
  ram[42015]  = 1;
  ram[42016]  = 1;
  ram[42017]  = 1;
  ram[42018]  = 1;
  ram[42019]  = 1;
  ram[42020]  = 1;
  ram[42021]  = 1;
  ram[42022]  = 1;
  ram[42023]  = 1;
  ram[42024]  = 1;
  ram[42025]  = 1;
  ram[42026]  = 1;
  ram[42027]  = 1;
  ram[42028]  = 1;
  ram[42029]  = 1;
  ram[42030]  = 1;
  ram[42031]  = 1;
  ram[42032]  = 1;
  ram[42033]  = 1;
  ram[42034]  = 1;
  ram[42035]  = 1;
  ram[42036]  = 1;
  ram[42037]  = 1;
  ram[42038]  = 1;
  ram[42039]  = 1;
  ram[42040]  = 1;
  ram[42041]  = 1;
  ram[42042]  = 1;
  ram[42043]  = 1;
  ram[42044]  = 1;
  ram[42045]  = 1;
  ram[42046]  = 1;
  ram[42047]  = 1;
  ram[42048]  = 1;
  ram[42049]  = 1;
  ram[42050]  = 1;
  ram[42051]  = 1;
  ram[42052]  = 1;
  ram[42053]  = 1;
  ram[42054]  = 1;
  ram[42055]  = 1;
  ram[42056]  = 1;
  ram[42057]  = 1;
  ram[42058]  = 1;
  ram[42059]  = 1;
  ram[42060]  = 1;
  ram[42061]  = 1;
  ram[42062]  = 1;
  ram[42063]  = 1;
  ram[42064]  = 1;
  ram[42065]  = 1;
  ram[42066]  = 1;
  ram[42067]  = 1;
  ram[42068]  = 1;
  ram[42069]  = 1;
  ram[42070]  = 1;
  ram[42071]  = 1;
  ram[42072]  = 1;
  ram[42073]  = 1;
  ram[42074]  = 1;
  ram[42075]  = 1;
  ram[42076]  = 1;
  ram[42077]  = 1;
  ram[42078]  = 1;
  ram[42079]  = 1;
  ram[42080]  = 1;
  ram[42081]  = 1;
  ram[42082]  = 1;
  ram[42083]  = 1;
  ram[42084]  = 1;
  ram[42085]  = 1;
  ram[42086]  = 1;
  ram[42087]  = 1;
  ram[42088]  = 1;
  ram[42089]  = 1;
  ram[42090]  = 1;
  ram[42091]  = 1;
  ram[42092]  = 1;
  ram[42093]  = 1;
  ram[42094]  = 1;
  ram[42095]  = 1;
  ram[42096]  = 1;
  ram[42097]  = 1;
  ram[42098]  = 1;
  ram[42099]  = 1;
  ram[42100]  = 1;
  ram[42101]  = 1;
  ram[42102]  = 1;
  ram[42103]  = 1;
  ram[42104]  = 1;
  ram[42105]  = 1;
  ram[42106]  = 1;
  ram[42107]  = 1;
  ram[42108]  = 1;
  ram[42109]  = 1;
  ram[42110]  = 1;
  ram[42111]  = 1;
  ram[42112]  = 1;
  ram[42113]  = 1;
  ram[42114]  = 1;
  ram[42115]  = 1;
  ram[42116]  = 1;
  ram[42117]  = 1;
  ram[42118]  = 1;
  ram[42119]  = 1;
  ram[42120]  = 1;
  ram[42121]  = 1;
  ram[42122]  = 1;
  ram[42123]  = 1;
  ram[42124]  = 1;
  ram[42125]  = 1;
  ram[42126]  = 1;
  ram[42127]  = 1;
  ram[42128]  = 1;
  ram[42129]  = 1;
  ram[42130]  = 1;
  ram[42131]  = 1;
  ram[42132]  = 1;
  ram[42133]  = 1;
  ram[42134]  = 1;
  ram[42135]  = 1;
  ram[42136]  = 1;
  ram[42137]  = 1;
  ram[42138]  = 1;
  ram[42139]  = 1;
  ram[42140]  = 1;
  ram[42141]  = 1;
  ram[42142]  = 1;
  ram[42143]  = 1;
  ram[42144]  = 1;
  ram[42145]  = 1;
  ram[42146]  = 1;
  ram[42147]  = 1;
  ram[42148]  = 1;
  ram[42149]  = 1;
  ram[42150]  = 1;
  ram[42151]  = 1;
  ram[42152]  = 1;
  ram[42153]  = 1;
  ram[42154]  = 1;
  ram[42155]  = 1;
  ram[42156]  = 1;
  ram[42157]  = 1;
  ram[42158]  = 1;
  ram[42159]  = 1;
  ram[42160]  = 1;
  ram[42161]  = 1;
  ram[42162]  = 1;
  ram[42163]  = 1;
  ram[42164]  = 1;
  ram[42165]  = 1;
  ram[42166]  = 1;
  ram[42167]  = 1;
  ram[42168]  = 1;
  ram[42169]  = 1;
  ram[42170]  = 1;
  ram[42171]  = 1;
  ram[42172]  = 1;
  ram[42173]  = 1;
  ram[42174]  = 1;
  ram[42175]  = 1;
  ram[42176]  = 1;
  ram[42177]  = 1;
  ram[42178]  = 1;
  ram[42179]  = 1;
  ram[42180]  = 1;
  ram[42181]  = 1;
  ram[42182]  = 1;
  ram[42183]  = 1;
  ram[42184]  = 1;
  ram[42185]  = 1;
  ram[42186]  = 1;
  ram[42187]  = 1;
  ram[42188]  = 1;
  ram[42189]  = 1;
  ram[42190]  = 1;
  ram[42191]  = 1;
  ram[42192]  = 1;
  ram[42193]  = 1;
  ram[42194]  = 1;
  ram[42195]  = 1;
  ram[42196]  = 1;
  ram[42197]  = 1;
  ram[42198]  = 1;
  ram[42199]  = 1;
  ram[42200]  = 1;
  ram[42201]  = 1;
  ram[42202]  = 1;
  ram[42203]  = 1;
  ram[42204]  = 1;
  ram[42205]  = 1;
  ram[42206]  = 1;
  ram[42207]  = 1;
  ram[42208]  = 1;
  ram[42209]  = 1;
  ram[42210]  = 1;
  ram[42211]  = 1;
  ram[42212]  = 1;
  ram[42213]  = 1;
  ram[42214]  = 1;
  ram[42215]  = 1;
  ram[42216]  = 1;
  ram[42217]  = 1;
  ram[42218]  = 1;
  ram[42219]  = 1;
  ram[42220]  = 1;
  ram[42221]  = 1;
  ram[42222]  = 1;
  ram[42223]  = 1;
  ram[42224]  = 1;
  ram[42225]  = 1;
  ram[42226]  = 1;
  ram[42227]  = 1;
  ram[42228]  = 1;
  ram[42229]  = 1;
  ram[42230]  = 1;
  ram[42231]  = 1;
  ram[42232]  = 1;
  ram[42233]  = 1;
  ram[42234]  = 1;
  ram[42235]  = 1;
  ram[42236]  = 1;
  ram[42237]  = 1;
  ram[42238]  = 1;
  ram[42239]  = 1;
  ram[42240]  = 1;
  ram[42241]  = 1;
  ram[42242]  = 1;
  ram[42243]  = 1;
  ram[42244]  = 1;
  ram[42245]  = 1;
  ram[42246]  = 1;
  ram[42247]  = 1;
  ram[42248]  = 1;
  ram[42249]  = 1;
  ram[42250]  = 1;
  ram[42251]  = 1;
  ram[42252]  = 1;
  ram[42253]  = 1;
  ram[42254]  = 1;
  ram[42255]  = 1;
  ram[42256]  = 1;
  ram[42257]  = 1;
  ram[42258]  = 1;
  ram[42259]  = 1;
  ram[42260]  = 1;
  ram[42261]  = 1;
  ram[42262]  = 1;
  ram[42263]  = 1;
  ram[42264]  = 1;
  ram[42265]  = 1;
  ram[42266]  = 1;
  ram[42267]  = 1;
  ram[42268]  = 1;
  ram[42269]  = 1;
  ram[42270]  = 1;
  ram[42271]  = 1;
  ram[42272]  = 1;
  ram[42273]  = 1;
  ram[42274]  = 1;
  ram[42275]  = 1;
  ram[42276]  = 1;
  ram[42277]  = 1;
  ram[42278]  = 1;
  ram[42279]  = 1;
  ram[42280]  = 1;
  ram[42281]  = 1;
  ram[42282]  = 1;
  ram[42283]  = 1;
  ram[42284]  = 1;
  ram[42285]  = 1;
  ram[42286]  = 1;
  ram[42287]  = 1;
  ram[42288]  = 1;
  ram[42289]  = 1;
  ram[42290]  = 1;
  ram[42291]  = 1;
  ram[42292]  = 1;
  ram[42293]  = 1;
  ram[42294]  = 1;
  ram[42295]  = 1;
  ram[42296]  = 1;
  ram[42297]  = 1;
  ram[42298]  = 1;
  ram[42299]  = 1;
  ram[42300]  = 1;
  ram[42301]  = 1;
  ram[42302]  = 1;
  ram[42303]  = 1;
  ram[42304]  = 1;
  ram[42305]  = 1;
  ram[42306]  = 1;
  ram[42307]  = 1;
  ram[42308]  = 1;
  ram[42309]  = 1;
  ram[42310]  = 1;
  ram[42311]  = 1;
  ram[42312]  = 1;
  ram[42313]  = 1;
  ram[42314]  = 1;
  ram[42315]  = 1;
  ram[42316]  = 1;
  ram[42317]  = 1;
  ram[42318]  = 1;
  ram[42319]  = 1;
  ram[42320]  = 1;
  ram[42321]  = 1;
  ram[42322]  = 1;
  ram[42323]  = 1;
  ram[42324]  = 1;
  ram[42325]  = 1;
  ram[42326]  = 1;
  ram[42327]  = 1;
  ram[42328]  = 1;
  ram[42329]  = 1;
  ram[42330]  = 1;
  ram[42331]  = 1;
  ram[42332]  = 1;
  ram[42333]  = 1;
  ram[42334]  = 1;
  ram[42335]  = 1;
  ram[42336]  = 1;
  ram[42337]  = 1;
  ram[42338]  = 1;
  ram[42339]  = 1;
  ram[42340]  = 1;
  ram[42341]  = 1;
  ram[42342]  = 1;
  ram[42343]  = 1;
  ram[42344]  = 1;
  ram[42345]  = 1;
  ram[42346]  = 1;
  ram[42347]  = 1;
  ram[42348]  = 1;
  ram[42349]  = 1;
  ram[42350]  = 1;
  ram[42351]  = 1;
  ram[42352]  = 1;
  ram[42353]  = 1;
  ram[42354]  = 1;
  ram[42355]  = 1;
  ram[42356]  = 1;
  ram[42357]  = 1;
  ram[42358]  = 1;
  ram[42359]  = 1;
  ram[42360]  = 1;
  ram[42361]  = 1;
  ram[42362]  = 1;
  ram[42363]  = 1;
  ram[42364]  = 1;
  ram[42365]  = 1;
  ram[42366]  = 1;
  ram[42367]  = 1;
  ram[42368]  = 1;
  ram[42369]  = 1;
  ram[42370]  = 1;
  ram[42371]  = 1;
  ram[42372]  = 1;
  ram[42373]  = 1;
  ram[42374]  = 1;
  ram[42375]  = 1;
  ram[42376]  = 1;
  ram[42377]  = 1;
  ram[42378]  = 1;
  ram[42379]  = 1;
  ram[42380]  = 1;
  ram[42381]  = 1;
  ram[42382]  = 1;
  ram[42383]  = 1;
  ram[42384]  = 1;
  ram[42385]  = 1;
  ram[42386]  = 1;
  ram[42387]  = 1;
  ram[42388]  = 1;
  ram[42389]  = 1;
  ram[42390]  = 1;
  ram[42391]  = 1;
  ram[42392]  = 1;
  ram[42393]  = 1;
  ram[42394]  = 1;
  ram[42395]  = 1;
  ram[42396]  = 1;
  ram[42397]  = 1;
  ram[42398]  = 1;
  ram[42399]  = 1;
  ram[42400]  = 1;
  ram[42401]  = 1;
  ram[42402]  = 1;
  ram[42403]  = 1;
  ram[42404]  = 1;
  ram[42405]  = 1;
  ram[42406]  = 1;
  ram[42407]  = 1;
  ram[42408]  = 1;
  ram[42409]  = 1;
  ram[42410]  = 1;
  ram[42411]  = 1;
  ram[42412]  = 1;
  ram[42413]  = 1;
  ram[42414]  = 1;
  ram[42415]  = 1;
  ram[42416]  = 1;
  ram[42417]  = 1;
  ram[42418]  = 1;
  ram[42419]  = 1;
  ram[42420]  = 1;
  ram[42421]  = 1;
  ram[42422]  = 1;
  ram[42423]  = 1;
  ram[42424]  = 1;
  ram[42425]  = 1;
  ram[42426]  = 1;
  ram[42427]  = 1;
  ram[42428]  = 1;
  ram[42429]  = 1;
  ram[42430]  = 1;
  ram[42431]  = 1;
  ram[42432]  = 1;
  ram[42433]  = 1;
  ram[42434]  = 1;
  ram[42435]  = 1;
  ram[42436]  = 1;
  ram[42437]  = 1;
  ram[42438]  = 1;
  ram[42439]  = 1;
  ram[42440]  = 1;
  ram[42441]  = 1;
  ram[42442]  = 1;
  ram[42443]  = 1;
  ram[42444]  = 1;
  ram[42445]  = 1;
  ram[42446]  = 1;
  ram[42447]  = 1;
  ram[42448]  = 1;
  ram[42449]  = 1;
  ram[42450]  = 1;
  ram[42451]  = 1;
  ram[42452]  = 1;
  ram[42453]  = 1;
  ram[42454]  = 1;
  ram[42455]  = 1;
  ram[42456]  = 1;
  ram[42457]  = 1;
  ram[42458]  = 1;
  ram[42459]  = 1;
  ram[42460]  = 1;
  ram[42461]  = 1;
  ram[42462]  = 1;
  ram[42463]  = 1;
  ram[42464]  = 1;
  ram[42465]  = 1;
  ram[42466]  = 1;
  ram[42467]  = 1;
  ram[42468]  = 1;
  ram[42469]  = 1;
  ram[42470]  = 1;
  ram[42471]  = 1;
  ram[42472]  = 1;
  ram[42473]  = 1;
  ram[42474]  = 1;
  ram[42475]  = 1;
  ram[42476]  = 1;
  ram[42477]  = 1;
  ram[42478]  = 1;
  ram[42479]  = 1;
  ram[42480]  = 1;
  ram[42481]  = 1;
  ram[42482]  = 1;
  ram[42483]  = 1;
  ram[42484]  = 1;
  ram[42485]  = 1;
  ram[42486]  = 1;
  ram[42487]  = 1;
  ram[42488]  = 1;
  ram[42489]  = 1;
  ram[42490]  = 1;
  ram[42491]  = 1;
  ram[42492]  = 1;
  ram[42493]  = 1;
  ram[42494]  = 1;
  ram[42495]  = 1;
  ram[42496]  = 1;
  ram[42497]  = 1;
  ram[42498]  = 1;
  ram[42499]  = 1;
  ram[42500]  = 1;
  ram[42501]  = 1;
  ram[42502]  = 1;
  ram[42503]  = 1;
  ram[42504]  = 1;
  ram[42505]  = 1;
  ram[42506]  = 1;
  ram[42507]  = 1;
  ram[42508]  = 1;
  ram[42509]  = 1;
  ram[42510]  = 1;
  ram[42511]  = 1;
  ram[42512]  = 1;
  ram[42513]  = 1;
  ram[42514]  = 1;
  ram[42515]  = 1;
  ram[42516]  = 1;
  ram[42517]  = 1;
  ram[42518]  = 1;
  ram[42519]  = 1;
  ram[42520]  = 1;
  ram[42521]  = 1;
  ram[42522]  = 1;
  ram[42523]  = 1;
  ram[42524]  = 1;
  ram[42525]  = 1;
  ram[42526]  = 1;
  ram[42527]  = 1;
  ram[42528]  = 1;
  ram[42529]  = 1;
  ram[42530]  = 1;
  ram[42531]  = 1;
  ram[42532]  = 1;
  ram[42533]  = 1;
  ram[42534]  = 1;
  ram[42535]  = 1;
  ram[42536]  = 1;
  ram[42537]  = 1;
  ram[42538]  = 1;
  ram[42539]  = 1;
  ram[42540]  = 1;
  ram[42541]  = 1;
  ram[42542]  = 1;
  ram[42543]  = 1;
  ram[42544]  = 1;
  ram[42545]  = 1;
  ram[42546]  = 1;
  ram[42547]  = 1;
  ram[42548]  = 1;
  ram[42549]  = 1;
  ram[42550]  = 1;
  ram[42551]  = 1;
  ram[42552]  = 1;
  ram[42553]  = 1;
  ram[42554]  = 1;
  ram[42555]  = 1;
  ram[42556]  = 1;
  ram[42557]  = 1;
  ram[42558]  = 1;
  ram[42559]  = 1;
  ram[42560]  = 1;
  ram[42561]  = 1;
  ram[42562]  = 1;
  ram[42563]  = 1;
  ram[42564]  = 1;
  ram[42565]  = 1;
  ram[42566]  = 1;
  ram[42567]  = 1;
  ram[42568]  = 1;
  ram[42569]  = 1;
  ram[42570]  = 1;
  ram[42571]  = 1;
  ram[42572]  = 1;
  ram[42573]  = 1;
  ram[42574]  = 1;
  ram[42575]  = 1;
  ram[42576]  = 1;
  ram[42577]  = 1;
  ram[42578]  = 1;
  ram[42579]  = 1;
  ram[42580]  = 1;
  ram[42581]  = 1;
  ram[42582]  = 1;
  ram[42583]  = 1;
  ram[42584]  = 1;
  ram[42585]  = 1;
  ram[42586]  = 1;
  ram[42587]  = 1;
  ram[42588]  = 1;
  ram[42589]  = 1;
  ram[42590]  = 1;
  ram[42591]  = 1;
  ram[42592]  = 1;
  ram[42593]  = 1;
  ram[42594]  = 1;
  ram[42595]  = 1;
  ram[42596]  = 1;
  ram[42597]  = 1;
  ram[42598]  = 1;
  ram[42599]  = 1;
  ram[42600]  = 1;
  ram[42601]  = 1;
  ram[42602]  = 1;
  ram[42603]  = 1;
  ram[42604]  = 1;
  ram[42605]  = 1;
  ram[42606]  = 1;
  ram[42607]  = 1;
  ram[42608]  = 1;
  ram[42609]  = 1;
  ram[42610]  = 1;
  ram[42611]  = 1;
  ram[42612]  = 1;
  ram[42613]  = 1;
  ram[42614]  = 1;
  ram[42615]  = 1;
  ram[42616]  = 1;
  ram[42617]  = 1;
  ram[42618]  = 1;
  ram[42619]  = 1;
  ram[42620]  = 1;
  ram[42621]  = 1;
  ram[42622]  = 1;
  ram[42623]  = 1;
  ram[42624]  = 1;
  ram[42625]  = 1;
  ram[42626]  = 1;
  ram[42627]  = 1;
  ram[42628]  = 1;
  ram[42629]  = 1;
  ram[42630]  = 1;
  ram[42631]  = 1;
  ram[42632]  = 1;
  ram[42633]  = 1;
  ram[42634]  = 1;
  ram[42635]  = 1;
  ram[42636]  = 1;
  ram[42637]  = 1;
  ram[42638]  = 1;
  ram[42639]  = 1;
  ram[42640]  = 1;
  ram[42641]  = 1;
  ram[42642]  = 1;
  ram[42643]  = 1;
  ram[42644]  = 1;
  ram[42645]  = 1;
  ram[42646]  = 1;
  ram[42647]  = 1;
  ram[42648]  = 1;
  ram[42649]  = 1;
  ram[42650]  = 1;
  ram[42651]  = 1;
  ram[42652]  = 1;
  ram[42653]  = 1;
  ram[42654]  = 1;
  ram[42655]  = 1;
  ram[42656]  = 1;
  ram[42657]  = 1;
  ram[42658]  = 1;
  ram[42659]  = 1;
  ram[42660]  = 1;
  ram[42661]  = 1;
  ram[42662]  = 1;
  ram[42663]  = 1;
  ram[42664]  = 1;
  ram[42665]  = 1;
  ram[42666]  = 1;
  ram[42667]  = 1;
  ram[42668]  = 1;
  ram[42669]  = 1;
  ram[42670]  = 1;
  ram[42671]  = 1;
  ram[42672]  = 1;
  ram[42673]  = 1;
  ram[42674]  = 1;
  ram[42675]  = 1;
  ram[42676]  = 1;
  ram[42677]  = 1;
  ram[42678]  = 1;
  ram[42679]  = 1;
  ram[42680]  = 1;
  ram[42681]  = 1;
  ram[42682]  = 1;
  ram[42683]  = 1;
  ram[42684]  = 1;
  ram[42685]  = 1;
  ram[42686]  = 1;
  ram[42687]  = 1;
  ram[42688]  = 1;
  ram[42689]  = 1;
  ram[42690]  = 1;
  ram[42691]  = 1;
  ram[42692]  = 1;
  ram[42693]  = 1;
  ram[42694]  = 1;
  ram[42695]  = 1;
  ram[42696]  = 1;
  ram[42697]  = 1;
  ram[42698]  = 1;
  ram[42699]  = 1;
  ram[42700]  = 1;
  ram[42701]  = 1;
  ram[42702]  = 1;
  ram[42703]  = 1;
  ram[42704]  = 1;
  ram[42705]  = 1;
  ram[42706]  = 1;
  ram[42707]  = 1;
  ram[42708]  = 1;
  ram[42709]  = 1;
  ram[42710]  = 1;
  ram[42711]  = 1;
  ram[42712]  = 1;
  ram[42713]  = 1;
  ram[42714]  = 1;
  ram[42715]  = 1;
  ram[42716]  = 1;
  ram[42717]  = 1;
  ram[42718]  = 1;
  ram[42719]  = 1;
  ram[42720]  = 1;
  ram[42721]  = 1;
  ram[42722]  = 1;
  ram[42723]  = 1;
  ram[42724]  = 1;
  ram[42725]  = 1;
  ram[42726]  = 1;
  ram[42727]  = 1;
  ram[42728]  = 1;
  ram[42729]  = 1;
  ram[42730]  = 1;
  ram[42731]  = 1;
  ram[42732]  = 1;
  ram[42733]  = 1;
  ram[42734]  = 1;
  ram[42735]  = 1;
  ram[42736]  = 1;
  ram[42737]  = 1;
  ram[42738]  = 1;
  ram[42739]  = 1;
  ram[42740]  = 1;
  ram[42741]  = 1;
  ram[42742]  = 1;
  ram[42743]  = 1;
  ram[42744]  = 1;
  ram[42745]  = 1;
  ram[42746]  = 1;
  ram[42747]  = 1;
  ram[42748]  = 1;
  ram[42749]  = 1;
  ram[42750]  = 1;
  ram[42751]  = 1;
  ram[42752]  = 1;
  ram[42753]  = 1;
  ram[42754]  = 1;
  ram[42755]  = 1;
  ram[42756]  = 1;
  ram[42757]  = 1;
  ram[42758]  = 1;
  ram[42759]  = 1;
  ram[42760]  = 1;
  ram[42761]  = 1;
  ram[42762]  = 1;
  ram[42763]  = 1;
  ram[42764]  = 1;
  ram[42765]  = 1;
  ram[42766]  = 1;
  ram[42767]  = 1;
  ram[42768]  = 1;
  ram[42769]  = 1;
  ram[42770]  = 1;
  ram[42771]  = 1;
  ram[42772]  = 1;
  ram[42773]  = 1;
  ram[42774]  = 1;
  ram[42775]  = 1;
  ram[42776]  = 1;
  ram[42777]  = 1;
  ram[42778]  = 1;
  ram[42779]  = 1;
  ram[42780]  = 1;
  ram[42781]  = 1;
  ram[42782]  = 1;
  ram[42783]  = 1;
  ram[42784]  = 1;
  ram[42785]  = 1;
  ram[42786]  = 1;
  ram[42787]  = 1;
  ram[42788]  = 1;
  ram[42789]  = 1;
  ram[42790]  = 1;
  ram[42791]  = 1;
  ram[42792]  = 1;
  ram[42793]  = 1;
  ram[42794]  = 1;
  ram[42795]  = 1;
  ram[42796]  = 1;
  ram[42797]  = 1;
  ram[42798]  = 1;
  ram[42799]  = 1;
  ram[42800]  = 1;
  ram[42801]  = 1;
  ram[42802]  = 1;
  ram[42803]  = 1;
  ram[42804]  = 1;
  ram[42805]  = 1;
  ram[42806]  = 1;
  ram[42807]  = 1;
  ram[42808]  = 1;
  ram[42809]  = 1;
  ram[42810]  = 1;
  ram[42811]  = 1;
  ram[42812]  = 1;
  ram[42813]  = 1;
  ram[42814]  = 1;
  ram[42815]  = 1;
  ram[42816]  = 1;
  ram[42817]  = 1;
  ram[42818]  = 1;
  ram[42819]  = 1;
  ram[42820]  = 1;
  ram[42821]  = 1;
  ram[42822]  = 1;
  ram[42823]  = 1;
  ram[42824]  = 1;
  ram[42825]  = 1;
  ram[42826]  = 1;
  ram[42827]  = 1;
  ram[42828]  = 1;
  ram[42829]  = 1;
  ram[42830]  = 1;
  ram[42831]  = 1;
  ram[42832]  = 1;
  ram[42833]  = 1;
  ram[42834]  = 1;
  ram[42835]  = 1;
  ram[42836]  = 1;
  ram[42837]  = 1;
  ram[42838]  = 1;
  ram[42839]  = 1;
  ram[42840]  = 1;
  ram[42841]  = 1;
  ram[42842]  = 1;
  ram[42843]  = 1;
  ram[42844]  = 1;
  ram[42845]  = 1;
  ram[42846]  = 1;
  ram[42847]  = 1;
  ram[42848]  = 1;
  ram[42849]  = 1;
  ram[42850]  = 1;
  ram[42851]  = 1;
  ram[42852]  = 1;
  ram[42853]  = 1;
  ram[42854]  = 1;
  ram[42855]  = 1;
  ram[42856]  = 1;
  ram[42857]  = 1;
  ram[42858]  = 1;
  ram[42859]  = 1;
  ram[42860]  = 1;
  ram[42861]  = 1;
  ram[42862]  = 1;
  ram[42863]  = 1;
  ram[42864]  = 1;
  ram[42865]  = 1;
  ram[42866]  = 1;
  ram[42867]  = 1;
  ram[42868]  = 1;
  ram[42869]  = 1;
  ram[42870]  = 1;
  ram[42871]  = 1;
  ram[42872]  = 1;
  ram[42873]  = 1;
  ram[42874]  = 1;
  ram[42875]  = 1;
  ram[42876]  = 1;
  ram[42877]  = 1;
  ram[42878]  = 1;
  ram[42879]  = 1;
  ram[42880]  = 1;
  ram[42881]  = 1;
  ram[42882]  = 1;
  ram[42883]  = 1;
  ram[42884]  = 1;
  ram[42885]  = 1;
  ram[42886]  = 1;
  ram[42887]  = 1;
  ram[42888]  = 1;
  ram[42889]  = 1;
  ram[42890]  = 1;
  ram[42891]  = 1;
  ram[42892]  = 1;
  ram[42893]  = 1;
  ram[42894]  = 1;
  ram[42895]  = 1;
  ram[42896]  = 1;
  ram[42897]  = 1;
  ram[42898]  = 1;
  ram[42899]  = 1;
  ram[42900]  = 1;
  ram[42901]  = 1;
  ram[42902]  = 1;
  ram[42903]  = 1;
  ram[42904]  = 1;
  ram[42905]  = 1;
  ram[42906]  = 1;
  ram[42907]  = 1;
  ram[42908]  = 1;
  ram[42909]  = 1;
  ram[42910]  = 1;
  ram[42911]  = 1;
  ram[42912]  = 1;
  ram[42913]  = 1;
  ram[42914]  = 1;
  ram[42915]  = 1;
  ram[42916]  = 1;
  ram[42917]  = 1;
  ram[42918]  = 1;
  ram[42919]  = 1;
  ram[42920]  = 1;
  ram[42921]  = 1;
  ram[42922]  = 1;
  ram[42923]  = 1;
  ram[42924]  = 1;
  ram[42925]  = 1;
  ram[42926]  = 1;
  ram[42927]  = 1;
  ram[42928]  = 1;
  ram[42929]  = 1;
  ram[42930]  = 1;
  ram[42931]  = 1;
  ram[42932]  = 1;
  ram[42933]  = 1;
  ram[42934]  = 1;
  ram[42935]  = 1;
  ram[42936]  = 1;
  ram[42937]  = 1;
  ram[42938]  = 1;
  ram[42939]  = 1;
  ram[42940]  = 1;
  ram[42941]  = 1;
  ram[42942]  = 1;
  ram[42943]  = 1;
  ram[42944]  = 1;
  ram[42945]  = 1;
  ram[42946]  = 1;
  ram[42947]  = 1;
  ram[42948]  = 1;
  ram[42949]  = 1;
  ram[42950]  = 1;
  ram[42951]  = 1;
  ram[42952]  = 1;
  ram[42953]  = 1;
  ram[42954]  = 1;
  ram[42955]  = 1;
  ram[42956]  = 1;
  ram[42957]  = 1;
  ram[42958]  = 1;
  ram[42959]  = 1;
  ram[42960]  = 1;
  ram[42961]  = 1;
  ram[42962]  = 1;
  ram[42963]  = 1;
  ram[42964]  = 1;
  ram[42965]  = 1;
  ram[42966]  = 1;
  ram[42967]  = 1;
  ram[42968]  = 1;
  ram[42969]  = 1;
  ram[42970]  = 1;
  ram[42971]  = 1;
  ram[42972]  = 1;
  ram[42973]  = 1;
  ram[42974]  = 1;
  ram[42975]  = 1;
  ram[42976]  = 1;
  ram[42977]  = 1;
  ram[42978]  = 1;
  ram[42979]  = 1;
  ram[42980]  = 1;
  ram[42981]  = 1;
  ram[42982]  = 1;
  ram[42983]  = 1;
  ram[42984]  = 1;
  ram[42985]  = 1;
  ram[42986]  = 1;
  ram[42987]  = 1;
  ram[42988]  = 1;
  ram[42989]  = 1;
  ram[42990]  = 1;
  ram[42991]  = 1;
  ram[42992]  = 1;
  ram[42993]  = 1;
  ram[42994]  = 1;
  ram[42995]  = 1;
  ram[42996]  = 1;
  ram[42997]  = 1;
  ram[42998]  = 1;
  ram[42999]  = 1;
  ram[43000]  = 1;
  ram[43001]  = 1;
  ram[43002]  = 1;
  ram[43003]  = 1;
  ram[43004]  = 1;
  ram[43005]  = 1;
  ram[43006]  = 1;
  ram[43007]  = 1;
  ram[43008]  = 1;
  ram[43009]  = 1;
  ram[43010]  = 1;
  ram[43011]  = 1;
  ram[43012]  = 1;
  ram[43013]  = 1;
  ram[43014]  = 1;
  ram[43015]  = 1;
  ram[43016]  = 1;
  ram[43017]  = 1;
  ram[43018]  = 1;
  ram[43019]  = 1;
  ram[43020]  = 1;
  ram[43021]  = 1;
  ram[43022]  = 1;
  ram[43023]  = 1;
  ram[43024]  = 1;
  ram[43025]  = 1;
  ram[43026]  = 1;
  ram[43027]  = 1;
  ram[43028]  = 1;
  ram[43029]  = 1;
  ram[43030]  = 1;
  ram[43031]  = 1;
  ram[43032]  = 1;
  ram[43033]  = 1;
  ram[43034]  = 1;
  ram[43035]  = 1;
  ram[43036]  = 1;
  ram[43037]  = 1;
  ram[43038]  = 1;
  ram[43039]  = 1;
  ram[43040]  = 1;
  ram[43041]  = 1;
  ram[43042]  = 1;
  ram[43043]  = 1;
  ram[43044]  = 1;
  ram[43045]  = 1;
  ram[43046]  = 1;
  ram[43047]  = 1;
  ram[43048]  = 1;
  ram[43049]  = 1;
  ram[43050]  = 1;
  ram[43051]  = 1;
  ram[43052]  = 1;
  ram[43053]  = 1;
  ram[43054]  = 1;
  ram[43055]  = 1;
  ram[43056]  = 1;
  ram[43057]  = 1;
  ram[43058]  = 1;
  ram[43059]  = 1;
  ram[43060]  = 1;
  ram[43061]  = 1;
  ram[43062]  = 1;
  ram[43063]  = 1;
  ram[43064]  = 1;
  ram[43065]  = 1;
  ram[43066]  = 1;
  ram[43067]  = 1;
  ram[43068]  = 1;
  ram[43069]  = 1;
  ram[43070]  = 1;
  ram[43071]  = 1;
  ram[43072]  = 1;
  ram[43073]  = 1;
  ram[43074]  = 1;
  ram[43075]  = 1;
  ram[43076]  = 1;
  ram[43077]  = 1;
  ram[43078]  = 1;
  ram[43079]  = 1;
  ram[43080]  = 1;
  ram[43081]  = 1;
  ram[43082]  = 1;
  ram[43083]  = 1;
  ram[43084]  = 1;
  ram[43085]  = 1;
  ram[43086]  = 1;
  ram[43087]  = 1;
  ram[43088]  = 1;
  ram[43089]  = 1;
  ram[43090]  = 1;
  ram[43091]  = 1;
  ram[43092]  = 1;
  ram[43093]  = 1;
  ram[43094]  = 1;
  ram[43095]  = 1;
  ram[43096]  = 1;
  ram[43097]  = 1;
  ram[43098]  = 1;
  ram[43099]  = 1;
  ram[43100]  = 1;
  ram[43101]  = 1;
  ram[43102]  = 1;
  ram[43103]  = 1;
  ram[43104]  = 1;
  ram[43105]  = 1;
  ram[43106]  = 1;
  ram[43107]  = 1;
  ram[43108]  = 1;
  ram[43109]  = 1;
  ram[43110]  = 1;
  ram[43111]  = 1;
  ram[43112]  = 1;
  ram[43113]  = 1;
  ram[43114]  = 1;
  ram[43115]  = 1;
  ram[43116]  = 1;
  ram[43117]  = 1;
  ram[43118]  = 1;
  ram[43119]  = 1;
  ram[43120]  = 1;
  ram[43121]  = 1;
  ram[43122]  = 1;
  ram[43123]  = 1;
  ram[43124]  = 1;
  ram[43125]  = 1;
  ram[43126]  = 1;
  ram[43127]  = 1;
  ram[43128]  = 1;
  ram[43129]  = 1;
  ram[43130]  = 1;
  ram[43131]  = 1;
  ram[43132]  = 1;
  ram[43133]  = 1;
  ram[43134]  = 1;
  ram[43135]  = 1;
  ram[43136]  = 1;
  ram[43137]  = 1;
  ram[43138]  = 1;
  ram[43139]  = 1;
  ram[43140]  = 1;
  ram[43141]  = 1;
  ram[43142]  = 1;
  ram[43143]  = 1;
  ram[43144]  = 1;
  ram[43145]  = 1;
  ram[43146]  = 1;
  ram[43147]  = 1;
  ram[43148]  = 1;
  ram[43149]  = 1;
  ram[43150]  = 1;
  ram[43151]  = 1;
  ram[43152]  = 1;
  ram[43153]  = 1;
  ram[43154]  = 1;
  ram[43155]  = 1;
  ram[43156]  = 1;
  ram[43157]  = 1;
  ram[43158]  = 1;
  ram[43159]  = 1;
  ram[43160]  = 1;
  ram[43161]  = 1;
  ram[43162]  = 1;
  ram[43163]  = 1;
  ram[43164]  = 1;
  ram[43165]  = 1;
  ram[43166]  = 1;
  ram[43167]  = 1;
  ram[43168]  = 1;
  ram[43169]  = 1;
  ram[43170]  = 1;
  ram[43171]  = 1;
  ram[43172]  = 1;
  ram[43173]  = 1;
  ram[43174]  = 1;
  ram[43175]  = 1;
  ram[43176]  = 1;
  ram[43177]  = 1;
  ram[43178]  = 1;
  ram[43179]  = 1;
  ram[43180]  = 1;
  ram[43181]  = 1;
  ram[43182]  = 1;
  ram[43183]  = 1;
  ram[43184]  = 1;
  ram[43185]  = 1;
  ram[43186]  = 1;
  ram[43187]  = 1;
  ram[43188]  = 1;
  ram[43189]  = 1;
  ram[43190]  = 1;
  ram[43191]  = 1;
  ram[43192]  = 1;
  ram[43193]  = 1;
  ram[43194]  = 1;
  ram[43195]  = 1;
  ram[43196]  = 1;
  ram[43197]  = 1;
  ram[43198]  = 1;
  ram[43199]  = 1;
  ram[43200]  = 1;
  ram[43201]  = 1;
  ram[43202]  = 1;
  ram[43203]  = 1;
  ram[43204]  = 1;
  ram[43205]  = 1;
  ram[43206]  = 1;
  ram[43207]  = 1;
  ram[43208]  = 1;
  ram[43209]  = 1;
  ram[43210]  = 1;
  ram[43211]  = 1;
  ram[43212]  = 1;
  ram[43213]  = 1;
  ram[43214]  = 1;
  ram[43215]  = 1;
  ram[43216]  = 1;
  ram[43217]  = 1;
  ram[43218]  = 1;
  ram[43219]  = 1;
  ram[43220]  = 1;
  ram[43221]  = 1;
  ram[43222]  = 1;
  ram[43223]  = 1;
  ram[43224]  = 1;
  ram[43225]  = 1;
  ram[43226]  = 1;
  ram[43227]  = 1;
  ram[43228]  = 1;
  ram[43229]  = 1;
  ram[43230]  = 1;
  ram[43231]  = 1;
  ram[43232]  = 1;
  ram[43233]  = 1;
  ram[43234]  = 1;
  ram[43235]  = 1;
  ram[43236]  = 1;
  ram[43237]  = 1;
  ram[43238]  = 1;
  ram[43239]  = 1;
  ram[43240]  = 1;
  ram[43241]  = 1;
  ram[43242]  = 1;
  ram[43243]  = 1;
  ram[43244]  = 1;
  ram[43245]  = 1;
  ram[43246]  = 1;
  ram[43247]  = 1;
  ram[43248]  = 1;
  ram[43249]  = 1;
  ram[43250]  = 1;
  ram[43251]  = 1;
  ram[43252]  = 1;
  ram[43253]  = 1;
  ram[43254]  = 1;
  ram[43255]  = 1;
  ram[43256]  = 1;
  ram[43257]  = 1;
  ram[43258]  = 1;
  ram[43259]  = 1;
  ram[43260]  = 1;
  ram[43261]  = 1;
  ram[43262]  = 1;
  ram[43263]  = 1;
  ram[43264]  = 1;
  ram[43265]  = 1;
  ram[43266]  = 1;
  ram[43267]  = 1;
  ram[43268]  = 1;
  ram[43269]  = 1;
  ram[43270]  = 1;
  ram[43271]  = 1;
  ram[43272]  = 1;
  ram[43273]  = 1;
  ram[43274]  = 1;
  ram[43275]  = 1;
  ram[43276]  = 1;
  ram[43277]  = 1;
  ram[43278]  = 1;
  ram[43279]  = 1;
  ram[43280]  = 1;
  ram[43281]  = 1;
  ram[43282]  = 1;
  ram[43283]  = 1;
  ram[43284]  = 1;
  ram[43285]  = 1;
  ram[43286]  = 1;
  ram[43287]  = 1;
  ram[43288]  = 1;
  ram[43289]  = 1;
  ram[43290]  = 1;
  ram[43291]  = 1;
  ram[43292]  = 1;
  ram[43293]  = 1;
  ram[43294]  = 1;
  ram[43295]  = 1;
  ram[43296]  = 1;
  ram[43297]  = 1;
  ram[43298]  = 1;
  ram[43299]  = 1;
  ram[43300]  = 1;
  ram[43301]  = 1;
  ram[43302]  = 1;
  ram[43303]  = 1;
  ram[43304]  = 1;
  ram[43305]  = 1;
  ram[43306]  = 1;
  ram[43307]  = 1;
  ram[43308]  = 1;
  ram[43309]  = 1;
  ram[43310]  = 1;
  ram[43311]  = 1;
  ram[43312]  = 1;
  ram[43313]  = 1;
  ram[43314]  = 1;
  ram[43315]  = 1;
  ram[43316]  = 1;
  ram[43317]  = 1;
  ram[43318]  = 1;
  ram[43319]  = 1;
  ram[43320]  = 1;
  ram[43321]  = 1;
  ram[43322]  = 1;
  ram[43323]  = 1;
  ram[43324]  = 1;
  ram[43325]  = 1;
  ram[43326]  = 1;
  ram[43327]  = 1;
  ram[43328]  = 1;
  ram[43329]  = 1;
  ram[43330]  = 1;
  ram[43331]  = 1;
  ram[43332]  = 1;
  ram[43333]  = 1;
  ram[43334]  = 1;
  ram[43335]  = 1;
  ram[43336]  = 1;
  ram[43337]  = 1;
  ram[43338]  = 1;
  ram[43339]  = 1;
  ram[43340]  = 1;
  ram[43341]  = 1;
  ram[43342]  = 1;
  ram[43343]  = 1;
  ram[43344]  = 1;
  ram[43345]  = 1;
  ram[43346]  = 1;
  ram[43347]  = 1;
  ram[43348]  = 1;
  ram[43349]  = 1;
  ram[43350]  = 1;
  ram[43351]  = 1;
  ram[43352]  = 1;
  ram[43353]  = 1;
  ram[43354]  = 1;
  ram[43355]  = 1;
  ram[43356]  = 1;
  ram[43357]  = 1;
  ram[43358]  = 1;
  ram[43359]  = 1;
  ram[43360]  = 1;
  ram[43361]  = 1;
  ram[43362]  = 1;
  ram[43363]  = 1;
  ram[43364]  = 1;
  ram[43365]  = 1;
  ram[43366]  = 1;
  ram[43367]  = 1;
  ram[43368]  = 1;
  ram[43369]  = 1;
  ram[43370]  = 1;
  ram[43371]  = 1;
  ram[43372]  = 1;
  ram[43373]  = 1;
  ram[43374]  = 1;
  ram[43375]  = 1;
  ram[43376]  = 1;
  ram[43377]  = 1;
  ram[43378]  = 1;
  ram[43379]  = 1;
  ram[43380]  = 1;
  ram[43381]  = 1;
  ram[43382]  = 1;
  ram[43383]  = 1;
  ram[43384]  = 1;
  ram[43385]  = 1;
  ram[43386]  = 1;
  ram[43387]  = 1;
  ram[43388]  = 1;
  ram[43389]  = 1;
  ram[43390]  = 1;
  ram[43391]  = 1;
  ram[43392]  = 1;
  ram[43393]  = 1;
  ram[43394]  = 1;
  ram[43395]  = 1;
  ram[43396]  = 1;
  ram[43397]  = 1;
  ram[43398]  = 1;
  ram[43399]  = 1;
  ram[43400]  = 1;
  ram[43401]  = 1;
  ram[43402]  = 1;
  ram[43403]  = 1;
  ram[43404]  = 1;
  ram[43405]  = 1;
  ram[43406]  = 1;
  ram[43407]  = 1;
  ram[43408]  = 1;
  ram[43409]  = 1;
  ram[43410]  = 1;
  ram[43411]  = 1;
  ram[43412]  = 1;
  ram[43413]  = 1;
  ram[43414]  = 1;
  ram[43415]  = 1;
  ram[43416]  = 1;
  ram[43417]  = 1;
  ram[43418]  = 1;
  ram[43419]  = 1;
  ram[43420]  = 1;
  ram[43421]  = 1;
  ram[43422]  = 1;
  ram[43423]  = 1;
  ram[43424]  = 1;
  ram[43425]  = 1;
  ram[43426]  = 1;
  ram[43427]  = 1;
  ram[43428]  = 1;
  ram[43429]  = 1;
  ram[43430]  = 1;
  ram[43431]  = 1;
  ram[43432]  = 1;
  ram[43433]  = 1;
  ram[43434]  = 1;
  ram[43435]  = 1;
  ram[43436]  = 1;
  ram[43437]  = 1;
  ram[43438]  = 1;
  ram[43439]  = 1;
  ram[43440]  = 1;
  ram[43441]  = 1;
  ram[43442]  = 1;
  ram[43443]  = 1;
  ram[43444]  = 1;
  ram[43445]  = 1;
  ram[43446]  = 1;
  ram[43447]  = 1;
  ram[43448]  = 1;
  ram[43449]  = 1;
  ram[43450]  = 1;
  ram[43451]  = 1;
  ram[43452]  = 1;
  ram[43453]  = 1;
  ram[43454]  = 1;
  ram[43455]  = 1;
  ram[43456]  = 1;
  ram[43457]  = 1;
  ram[43458]  = 1;
  ram[43459]  = 1;
  ram[43460]  = 1;
  ram[43461]  = 1;
  ram[43462]  = 1;
  ram[43463]  = 1;
  ram[43464]  = 1;
  ram[43465]  = 1;
  ram[43466]  = 1;
  ram[43467]  = 1;
  ram[43468]  = 1;
  ram[43469]  = 1;
  ram[43470]  = 1;
  ram[43471]  = 1;
  ram[43472]  = 1;
  ram[43473]  = 1;
  ram[43474]  = 1;
  ram[43475]  = 1;
  ram[43476]  = 1;
  ram[43477]  = 1;
  ram[43478]  = 1;
  ram[43479]  = 1;
  ram[43480]  = 1;
  ram[43481]  = 1;
  ram[43482]  = 1;
  ram[43483]  = 1;
  ram[43484]  = 1;
  ram[43485]  = 1;
  ram[43486]  = 1;
  ram[43487]  = 1;
  ram[43488]  = 1;
  ram[43489]  = 1;
  ram[43490]  = 1;
  ram[43491]  = 1;
  ram[43492]  = 1;
  ram[43493]  = 1;
  ram[43494]  = 1;
  ram[43495]  = 1;
  ram[43496]  = 1;
  ram[43497]  = 1;
  ram[43498]  = 1;
  ram[43499]  = 1;
  ram[43500]  = 1;
  ram[43501]  = 1;
  ram[43502]  = 1;
  ram[43503]  = 1;
  ram[43504]  = 1;
  ram[43505]  = 1;
  ram[43506]  = 1;
  ram[43507]  = 1;
  ram[43508]  = 1;
  ram[43509]  = 1;
  ram[43510]  = 1;
  ram[43511]  = 1;
  ram[43512]  = 1;
  ram[43513]  = 1;
  ram[43514]  = 1;
  ram[43515]  = 1;
  ram[43516]  = 1;
  ram[43517]  = 1;
  ram[43518]  = 1;
  ram[43519]  = 1;
  ram[43520]  = 1;
  ram[43521]  = 1;
  ram[43522]  = 1;
  ram[43523]  = 1;
  ram[43524]  = 1;
  ram[43525]  = 1;
  ram[43526]  = 1;
  ram[43527]  = 1;
  ram[43528]  = 1;
  ram[43529]  = 1;
  ram[43530]  = 1;
  ram[43531]  = 1;
  ram[43532]  = 1;
  ram[43533]  = 1;
  ram[43534]  = 1;
  ram[43535]  = 1;
  ram[43536]  = 1;
  ram[43537]  = 1;
  ram[43538]  = 1;
  ram[43539]  = 1;
  ram[43540]  = 1;
  ram[43541]  = 1;
  ram[43542]  = 1;
  ram[43543]  = 1;
  ram[43544]  = 1;
  ram[43545]  = 1;
  ram[43546]  = 1;
  ram[43547]  = 1;
  ram[43548]  = 1;
  ram[43549]  = 1;
  ram[43550]  = 1;
  ram[43551]  = 1;
  ram[43552]  = 1;
  ram[43553]  = 1;
  ram[43554]  = 1;
  ram[43555]  = 1;
  ram[43556]  = 1;
  ram[43557]  = 1;
  ram[43558]  = 1;
  ram[43559]  = 1;
  ram[43560]  = 1;
  ram[43561]  = 1;
  ram[43562]  = 1;
  ram[43563]  = 1;
  ram[43564]  = 1;
  ram[43565]  = 1;
  ram[43566]  = 1;
  ram[43567]  = 1;
  ram[43568]  = 1;
  ram[43569]  = 1;
  ram[43570]  = 1;
  ram[43571]  = 1;
  ram[43572]  = 1;
  ram[43573]  = 1;
  ram[43574]  = 1;
  ram[43575]  = 1;
  ram[43576]  = 1;
  ram[43577]  = 1;
  ram[43578]  = 1;
  ram[43579]  = 1;
  ram[43580]  = 1;
  ram[43581]  = 1;
  ram[43582]  = 1;
  ram[43583]  = 1;
  ram[43584]  = 1;
  ram[43585]  = 1;
  ram[43586]  = 1;
  ram[43587]  = 1;
  ram[43588]  = 1;
  ram[43589]  = 1;
  ram[43590]  = 1;
  ram[43591]  = 1;
  ram[43592]  = 1;
  ram[43593]  = 1;
  ram[43594]  = 1;
  ram[43595]  = 1;
  ram[43596]  = 1;
  ram[43597]  = 1;
  ram[43598]  = 1;
  ram[43599]  = 1;
  ram[43600]  = 1;
  ram[43601]  = 1;
  ram[43602]  = 1;
  ram[43603]  = 1;
  ram[43604]  = 1;
  ram[43605]  = 1;
  ram[43606]  = 1;
  ram[43607]  = 1;
  ram[43608]  = 1;
  ram[43609]  = 1;
  ram[43610]  = 1;
  ram[43611]  = 1;
  ram[43612]  = 1;
  ram[43613]  = 1;
  ram[43614]  = 1;
  ram[43615]  = 1;
  ram[43616]  = 1;
  ram[43617]  = 1;
  ram[43618]  = 1;
  ram[43619]  = 1;
  ram[43620]  = 1;
  ram[43621]  = 1;
  ram[43622]  = 1;
  ram[43623]  = 1;
  ram[43624]  = 1;
  ram[43625]  = 1;
  ram[43626]  = 1;
  ram[43627]  = 1;
  ram[43628]  = 1;
  ram[43629]  = 1;
  ram[43630]  = 1;
  ram[43631]  = 1;
  ram[43632]  = 1;
  ram[43633]  = 1;
  ram[43634]  = 1;
  ram[43635]  = 1;
  ram[43636]  = 1;
  ram[43637]  = 1;
  ram[43638]  = 1;
  ram[43639]  = 1;
  ram[43640]  = 1;
  ram[43641]  = 1;
  ram[43642]  = 1;
  ram[43643]  = 1;
  ram[43644]  = 1;
  ram[43645]  = 1;
  ram[43646]  = 1;
  ram[43647]  = 1;
  ram[43648]  = 1;
  ram[43649]  = 1;
  ram[43650]  = 1;
  ram[43651]  = 1;
  ram[43652]  = 1;
  ram[43653]  = 1;
  ram[43654]  = 1;
  ram[43655]  = 1;
  ram[43656]  = 1;
  ram[43657]  = 1;
  ram[43658]  = 1;
  ram[43659]  = 1;
  ram[43660]  = 1;
  ram[43661]  = 1;
  ram[43662]  = 1;
  ram[43663]  = 1;
  ram[43664]  = 1;
  ram[43665]  = 1;
  ram[43666]  = 1;
  ram[43667]  = 1;
  ram[43668]  = 1;
  ram[43669]  = 1;
  ram[43670]  = 1;
  ram[43671]  = 1;
  ram[43672]  = 1;
  ram[43673]  = 1;
  ram[43674]  = 1;
  ram[43675]  = 1;
  ram[43676]  = 1;
  ram[43677]  = 1;
  ram[43678]  = 1;
  ram[43679]  = 1;
  ram[43680]  = 1;
  ram[43681]  = 1;
  ram[43682]  = 1;
  ram[43683]  = 1;
  ram[43684]  = 1;
  ram[43685]  = 1;
  ram[43686]  = 1;
  ram[43687]  = 1;
  ram[43688]  = 1;
  ram[43689]  = 1;
  ram[43690]  = 1;
  ram[43691]  = 1;
  ram[43692]  = 1;
  ram[43693]  = 1;
  ram[43694]  = 1;
  ram[43695]  = 1;
  ram[43696]  = 1;
  ram[43697]  = 1;
  ram[43698]  = 1;
  ram[43699]  = 1;
  ram[43700]  = 1;
  ram[43701]  = 1;
  ram[43702]  = 1;
  ram[43703]  = 1;
  ram[43704]  = 1;
  ram[43705]  = 1;
  ram[43706]  = 1;
  ram[43707]  = 1;
  ram[43708]  = 1;
  ram[43709]  = 1;
  ram[43710]  = 1;
  ram[43711]  = 1;
  ram[43712]  = 1;
  ram[43713]  = 1;
  ram[43714]  = 1;
  ram[43715]  = 1;
  ram[43716]  = 1;
  ram[43717]  = 1;
  ram[43718]  = 1;
  ram[43719]  = 1;
  ram[43720]  = 1;
  ram[43721]  = 1;
  ram[43722]  = 1;
  ram[43723]  = 1;
  ram[43724]  = 1;
  ram[43725]  = 1;
  ram[43726]  = 1;
  ram[43727]  = 1;
  ram[43728]  = 1;
  ram[43729]  = 1;
  ram[43730]  = 1;
  ram[43731]  = 1;
  ram[43732]  = 1;
  ram[43733]  = 1;
  ram[43734]  = 1;
  ram[43735]  = 1;
  ram[43736]  = 1;
  ram[43737]  = 1;
  ram[43738]  = 1;
  ram[43739]  = 1;
  ram[43740]  = 1;
  ram[43741]  = 1;
  ram[43742]  = 1;
  ram[43743]  = 1;
  ram[43744]  = 1;
  ram[43745]  = 1;
  ram[43746]  = 1;
  ram[43747]  = 1;
  ram[43748]  = 1;
  ram[43749]  = 1;
  ram[43750]  = 1;
  ram[43751]  = 1;
  ram[43752]  = 1;
  ram[43753]  = 1;
  ram[43754]  = 1;
  ram[43755]  = 1;
  ram[43756]  = 1;
  ram[43757]  = 1;
  ram[43758]  = 1;
  ram[43759]  = 1;
  ram[43760]  = 1;
  ram[43761]  = 1;
  ram[43762]  = 1;
  ram[43763]  = 1;
  ram[43764]  = 1;
  ram[43765]  = 1;
  ram[43766]  = 1;
  ram[43767]  = 1;
  ram[43768]  = 1;
  ram[43769]  = 1;
  ram[43770]  = 1;
  ram[43771]  = 1;
  ram[43772]  = 1;
  ram[43773]  = 1;
  ram[43774]  = 1;
  ram[43775]  = 1;
  ram[43776]  = 1;
  ram[43777]  = 1;
  ram[43778]  = 1;
  ram[43779]  = 1;
  ram[43780]  = 1;
  ram[43781]  = 1;
  ram[43782]  = 1;
  ram[43783]  = 1;
  ram[43784]  = 1;
  ram[43785]  = 1;
  ram[43786]  = 1;
  ram[43787]  = 1;
  ram[43788]  = 1;
  ram[43789]  = 1;
  ram[43790]  = 1;
  ram[43791]  = 1;
  ram[43792]  = 1;
  ram[43793]  = 1;
  ram[43794]  = 1;
  ram[43795]  = 1;
  ram[43796]  = 1;
  ram[43797]  = 1;
  ram[43798]  = 1;
  ram[43799]  = 1;
  ram[43800]  = 1;
  ram[43801]  = 1;
  ram[43802]  = 1;
  ram[43803]  = 1;
  ram[43804]  = 1;
  ram[43805]  = 1;
  ram[43806]  = 1;
  ram[43807]  = 1;
  ram[43808]  = 1;
  ram[43809]  = 1;
  ram[43810]  = 1;
  ram[43811]  = 1;
  ram[43812]  = 1;
  ram[43813]  = 1;
  ram[43814]  = 1;
  ram[43815]  = 1;
  ram[43816]  = 1;
  ram[43817]  = 1;
  ram[43818]  = 1;
  ram[43819]  = 1;
  ram[43820]  = 1;
  ram[43821]  = 1;
  ram[43822]  = 1;
  ram[43823]  = 1;
  ram[43824]  = 1;
  ram[43825]  = 1;
  ram[43826]  = 1;
  ram[43827]  = 1;
  ram[43828]  = 1;
  ram[43829]  = 1;
  ram[43830]  = 1;
  ram[43831]  = 1;
  ram[43832]  = 1;
  ram[43833]  = 1;
  ram[43834]  = 1;
  ram[43835]  = 1;
  ram[43836]  = 1;
  ram[43837]  = 1;
  ram[43838]  = 1;
  ram[43839]  = 1;
  ram[43840]  = 1;
  ram[43841]  = 1;
  ram[43842]  = 1;
  ram[43843]  = 1;
  ram[43844]  = 1;
  ram[43845]  = 1;
  ram[43846]  = 1;
  ram[43847]  = 1;
  ram[43848]  = 1;
  ram[43849]  = 1;
  ram[43850]  = 1;
  ram[43851]  = 1;
  ram[43852]  = 1;
  ram[43853]  = 1;
  ram[43854]  = 1;
  ram[43855]  = 1;
  ram[43856]  = 1;
  ram[43857]  = 1;
  ram[43858]  = 1;
  ram[43859]  = 1;
  ram[43860]  = 1;
  ram[43861]  = 1;
  ram[43862]  = 1;
  ram[43863]  = 1;
  ram[43864]  = 1;
  ram[43865]  = 1;
  ram[43866]  = 1;
  ram[43867]  = 1;
  ram[43868]  = 1;
  ram[43869]  = 1;
  ram[43870]  = 1;
  ram[43871]  = 1;
  ram[43872]  = 1;
  ram[43873]  = 1;
  ram[43874]  = 1;
  ram[43875]  = 1;
  ram[43876]  = 1;
  ram[43877]  = 1;
  ram[43878]  = 1;
  ram[43879]  = 1;
  ram[43880]  = 1;
  ram[43881]  = 1;
  ram[43882]  = 1;
  ram[43883]  = 1;
  ram[43884]  = 1;
  ram[43885]  = 1;
  ram[43886]  = 1;
  ram[43887]  = 1;
  ram[43888]  = 1;
  ram[43889]  = 1;
  ram[43890]  = 1;
  ram[43891]  = 1;
  ram[43892]  = 1;
  ram[43893]  = 1;
  ram[43894]  = 1;
  ram[43895]  = 1;
  ram[43896]  = 1;
  ram[43897]  = 1;
  ram[43898]  = 1;
  ram[43899]  = 1;
  ram[43900]  = 1;
  ram[43901]  = 1;
  ram[43902]  = 1;
  ram[43903]  = 1;
  ram[43904]  = 1;
  ram[43905]  = 1;
  ram[43906]  = 1;
  ram[43907]  = 1;
  ram[43908]  = 1;
  ram[43909]  = 1;
  ram[43910]  = 1;
  ram[43911]  = 1;
  ram[43912]  = 1;
  ram[43913]  = 1;
  ram[43914]  = 1;
  ram[43915]  = 1;
  ram[43916]  = 1;
  ram[43917]  = 1;
  ram[43918]  = 1;
  ram[43919]  = 1;
  ram[43920]  = 1;
  ram[43921]  = 1;
  ram[43922]  = 1;
  ram[43923]  = 1;
  ram[43924]  = 1;
  ram[43925]  = 1;
  ram[43926]  = 1;
  ram[43927]  = 1;
  ram[43928]  = 1;
  ram[43929]  = 1;
  ram[43930]  = 1;
  ram[43931]  = 1;
  ram[43932]  = 1;
  ram[43933]  = 1;
  ram[43934]  = 1;
  ram[43935]  = 1;
  ram[43936]  = 1;
  ram[43937]  = 1;
  ram[43938]  = 1;
  ram[43939]  = 1;
  ram[43940]  = 1;
  ram[43941]  = 1;
  ram[43942]  = 1;
  ram[43943]  = 1;
  ram[43944]  = 1;
  ram[43945]  = 1;
  ram[43946]  = 1;
  ram[43947]  = 1;
  ram[43948]  = 1;
  ram[43949]  = 1;
  ram[43950]  = 1;
  ram[43951]  = 1;
  ram[43952]  = 1;
  ram[43953]  = 1;
  ram[43954]  = 1;
  ram[43955]  = 1;
  ram[43956]  = 1;
  ram[43957]  = 1;
  ram[43958]  = 1;
  ram[43959]  = 1;
  ram[43960]  = 1;
  ram[43961]  = 1;
  ram[43962]  = 1;
  ram[43963]  = 1;
  ram[43964]  = 1;
  ram[43965]  = 1;
  ram[43966]  = 1;
  ram[43967]  = 1;
  ram[43968]  = 1;
  ram[43969]  = 1;
  ram[43970]  = 1;
  ram[43971]  = 1;
  ram[43972]  = 1;
  ram[43973]  = 1;
  ram[43974]  = 1;
  ram[43975]  = 1;
  ram[43976]  = 1;
  ram[43977]  = 1;
  ram[43978]  = 1;
  ram[43979]  = 1;
  ram[43980]  = 1;
  ram[43981]  = 1;
  ram[43982]  = 1;
  ram[43983]  = 1;
  ram[43984]  = 1;
  ram[43985]  = 1;
  ram[43986]  = 1;
  ram[43987]  = 1;
  ram[43988]  = 1;
  ram[43989]  = 1;
  ram[43990]  = 1;
  ram[43991]  = 1;
  ram[43992]  = 1;
  ram[43993]  = 1;
  ram[43994]  = 1;
  ram[43995]  = 1;
  ram[43996]  = 1;
  ram[43997]  = 1;
  ram[43998]  = 1;
  ram[43999]  = 1;
  ram[44000]  = 1;
  ram[44001]  = 1;
  ram[44002]  = 1;
  ram[44003]  = 1;
  ram[44004]  = 1;
  ram[44005]  = 1;
  ram[44006]  = 1;
  ram[44007]  = 1;
  ram[44008]  = 1;
  ram[44009]  = 1;
  ram[44010]  = 1;
  ram[44011]  = 1;
  ram[44012]  = 1;
  ram[44013]  = 1;
  ram[44014]  = 1;
  ram[44015]  = 1;
  ram[44016]  = 1;
  ram[44017]  = 1;
  ram[44018]  = 1;
  ram[44019]  = 1;
  ram[44020]  = 1;
  ram[44021]  = 1;
  ram[44022]  = 1;
  ram[44023]  = 1;
  ram[44024]  = 1;
  ram[44025]  = 1;
  ram[44026]  = 1;
  ram[44027]  = 1;
  ram[44028]  = 1;
  ram[44029]  = 1;
  ram[44030]  = 1;
  ram[44031]  = 1;
  ram[44032]  = 1;
  ram[44033]  = 1;
  ram[44034]  = 1;
  ram[44035]  = 1;
  ram[44036]  = 1;
  ram[44037]  = 1;
  ram[44038]  = 1;
  ram[44039]  = 1;
  ram[44040]  = 1;
  ram[44041]  = 1;
  ram[44042]  = 1;
  ram[44043]  = 1;
  ram[44044]  = 1;
  ram[44045]  = 1;
  ram[44046]  = 1;
  ram[44047]  = 1;
  ram[44048]  = 1;
  ram[44049]  = 1;
  ram[44050]  = 1;
  ram[44051]  = 1;
  ram[44052]  = 1;
  ram[44053]  = 1;
  ram[44054]  = 1;
  ram[44055]  = 1;
  ram[44056]  = 1;
  ram[44057]  = 1;
  ram[44058]  = 1;
  ram[44059]  = 1;
  ram[44060]  = 1;
  ram[44061]  = 1;
  ram[44062]  = 1;
  ram[44063]  = 1;
  ram[44064]  = 1;
  ram[44065]  = 1;
  ram[44066]  = 1;
  ram[44067]  = 1;
  ram[44068]  = 1;
  ram[44069]  = 1;
  ram[44070]  = 1;
  ram[44071]  = 1;
  ram[44072]  = 1;
  ram[44073]  = 1;
  ram[44074]  = 1;
  ram[44075]  = 1;
  ram[44076]  = 1;
  ram[44077]  = 1;
  ram[44078]  = 1;
  ram[44079]  = 1;
  ram[44080]  = 1;
  ram[44081]  = 1;
  ram[44082]  = 1;
  ram[44083]  = 1;
  ram[44084]  = 1;
  ram[44085]  = 1;
  ram[44086]  = 1;
  ram[44087]  = 1;
  ram[44088]  = 1;
  ram[44089]  = 1;
  ram[44090]  = 1;
  ram[44091]  = 1;
  ram[44092]  = 1;
  ram[44093]  = 1;
  ram[44094]  = 1;
  ram[44095]  = 1;
  ram[44096]  = 1;
  ram[44097]  = 1;
  ram[44098]  = 1;
  ram[44099]  = 1;
  ram[44100]  = 1;
  ram[44101]  = 1;
  ram[44102]  = 1;
  ram[44103]  = 1;
  ram[44104]  = 1;
  ram[44105]  = 1;
  ram[44106]  = 1;
  ram[44107]  = 1;
  ram[44108]  = 1;
  ram[44109]  = 1;
  ram[44110]  = 1;
  ram[44111]  = 1;
  ram[44112]  = 1;
  ram[44113]  = 1;
  ram[44114]  = 1;
  ram[44115]  = 1;
  ram[44116]  = 1;
  ram[44117]  = 1;
  ram[44118]  = 1;
  ram[44119]  = 1;
  ram[44120]  = 1;
  ram[44121]  = 1;
  ram[44122]  = 1;
  ram[44123]  = 1;
  ram[44124]  = 1;
  ram[44125]  = 1;
  ram[44126]  = 1;
  ram[44127]  = 1;
  ram[44128]  = 1;
  ram[44129]  = 1;
  ram[44130]  = 1;
  ram[44131]  = 1;
  ram[44132]  = 1;
  ram[44133]  = 1;
  ram[44134]  = 1;
  ram[44135]  = 1;
  ram[44136]  = 1;
  ram[44137]  = 1;
  ram[44138]  = 1;
  ram[44139]  = 1;
  ram[44140]  = 1;
  ram[44141]  = 1;
  ram[44142]  = 1;
  ram[44143]  = 1;
  ram[44144]  = 1;
  ram[44145]  = 1;
  ram[44146]  = 1;
  ram[44147]  = 1;
  ram[44148]  = 1;
  ram[44149]  = 1;
  ram[44150]  = 1;
  ram[44151]  = 1;
  ram[44152]  = 1;
  ram[44153]  = 1;
  ram[44154]  = 1;
  ram[44155]  = 1;
  ram[44156]  = 1;
  ram[44157]  = 1;
  ram[44158]  = 1;
  ram[44159]  = 1;
  ram[44160]  = 1;
  ram[44161]  = 1;
  ram[44162]  = 1;
  ram[44163]  = 1;
  ram[44164]  = 1;
  ram[44165]  = 1;
  ram[44166]  = 1;
  ram[44167]  = 1;
  ram[44168]  = 1;
  ram[44169]  = 1;
  ram[44170]  = 1;
  ram[44171]  = 1;
  ram[44172]  = 1;
  ram[44173]  = 1;
  ram[44174]  = 1;
  ram[44175]  = 1;
  ram[44176]  = 1;
  ram[44177]  = 1;
  ram[44178]  = 1;
  ram[44179]  = 1;
  ram[44180]  = 1;
  ram[44181]  = 1;
  ram[44182]  = 1;
  ram[44183]  = 1;
  ram[44184]  = 1;
  ram[44185]  = 1;
  ram[44186]  = 1;
  ram[44187]  = 1;
  ram[44188]  = 1;
  ram[44189]  = 1;
  ram[44190]  = 1;
  ram[44191]  = 1;
  ram[44192]  = 1;
  ram[44193]  = 1;
  ram[44194]  = 1;
  ram[44195]  = 1;
  ram[44196]  = 1;
  ram[44197]  = 1;
  ram[44198]  = 1;
  ram[44199]  = 1;
  ram[44200]  = 1;
  ram[44201]  = 1;
  ram[44202]  = 1;
  ram[44203]  = 1;
  ram[44204]  = 1;
  ram[44205]  = 1;
  ram[44206]  = 1;
  ram[44207]  = 1;
  ram[44208]  = 1;
  ram[44209]  = 1;
  ram[44210]  = 1;
  ram[44211]  = 1;
  ram[44212]  = 1;
  ram[44213]  = 1;
  ram[44214]  = 1;
  ram[44215]  = 1;
  ram[44216]  = 1;
  ram[44217]  = 1;
  ram[44218]  = 1;
  ram[44219]  = 1;
  ram[44220]  = 1;
  ram[44221]  = 1;
  ram[44222]  = 1;
  ram[44223]  = 1;
  ram[44224]  = 1;
  ram[44225]  = 1;
  ram[44226]  = 1;
  ram[44227]  = 1;
  ram[44228]  = 1;
  ram[44229]  = 1;
  ram[44230]  = 1;
  ram[44231]  = 1;
  ram[44232]  = 1;
  ram[44233]  = 1;
  ram[44234]  = 1;
  ram[44235]  = 1;
  ram[44236]  = 1;
  ram[44237]  = 1;
  ram[44238]  = 1;
  ram[44239]  = 1;
  ram[44240]  = 1;
  ram[44241]  = 1;
  ram[44242]  = 1;
  ram[44243]  = 1;
  ram[44244]  = 1;
  ram[44245]  = 1;
  ram[44246]  = 1;
  ram[44247]  = 1;
  ram[44248]  = 1;
  ram[44249]  = 1;
  ram[44250]  = 1;
  ram[44251]  = 1;
  ram[44252]  = 1;
  ram[44253]  = 1;
  ram[44254]  = 1;
  ram[44255]  = 1;
  ram[44256]  = 1;
  ram[44257]  = 1;
  ram[44258]  = 1;
  ram[44259]  = 1;
  ram[44260]  = 1;
  ram[44261]  = 1;
  ram[44262]  = 1;
  ram[44263]  = 1;
  ram[44264]  = 1;
  ram[44265]  = 1;
  ram[44266]  = 1;
  ram[44267]  = 1;
  ram[44268]  = 1;
  ram[44269]  = 1;
  ram[44270]  = 1;
  ram[44271]  = 1;
  ram[44272]  = 1;
  ram[44273]  = 1;
  ram[44274]  = 1;
  ram[44275]  = 1;
  ram[44276]  = 1;
  ram[44277]  = 1;
  ram[44278]  = 1;
  ram[44279]  = 1;
  ram[44280]  = 1;
  ram[44281]  = 1;
  ram[44282]  = 1;
  ram[44283]  = 1;
  ram[44284]  = 1;
  ram[44285]  = 1;
  ram[44286]  = 1;
  ram[44287]  = 1;
  ram[44288]  = 1;
  ram[44289]  = 1;
  ram[44290]  = 1;
  ram[44291]  = 1;
  ram[44292]  = 1;
  ram[44293]  = 1;
  ram[44294]  = 1;
  ram[44295]  = 1;
  ram[44296]  = 1;
  ram[44297]  = 1;
  ram[44298]  = 1;
  ram[44299]  = 1;
  ram[44300]  = 1;
  ram[44301]  = 1;
  ram[44302]  = 1;
  ram[44303]  = 1;
  ram[44304]  = 1;
  ram[44305]  = 1;
  ram[44306]  = 1;
  ram[44307]  = 1;
  ram[44308]  = 1;
  ram[44309]  = 1;
  ram[44310]  = 1;
  ram[44311]  = 1;
  ram[44312]  = 1;
  ram[44313]  = 1;
  ram[44314]  = 1;
  ram[44315]  = 1;
  ram[44316]  = 1;
  ram[44317]  = 1;
  ram[44318]  = 1;
  ram[44319]  = 1;
  ram[44320]  = 1;
  ram[44321]  = 1;
  ram[44322]  = 1;
  ram[44323]  = 1;
  ram[44324]  = 1;
  ram[44325]  = 1;
  ram[44326]  = 1;
  ram[44327]  = 1;
  ram[44328]  = 1;
  ram[44329]  = 1;
  ram[44330]  = 1;
  ram[44331]  = 1;
  ram[44332]  = 1;
  ram[44333]  = 1;
  ram[44334]  = 1;
  ram[44335]  = 1;
  ram[44336]  = 1;
  ram[44337]  = 1;
  ram[44338]  = 1;
  ram[44339]  = 1;
  ram[44340]  = 1;
  ram[44341]  = 1;
  ram[44342]  = 1;
  ram[44343]  = 1;
  ram[44344]  = 1;
  ram[44345]  = 1;
  ram[44346]  = 1;
  ram[44347]  = 1;
  ram[44348]  = 1;
  ram[44349]  = 1;
  ram[44350]  = 1;
  ram[44351]  = 1;
  ram[44352]  = 1;
  ram[44353]  = 1;
  ram[44354]  = 1;
  ram[44355]  = 1;
  ram[44356]  = 1;
  ram[44357]  = 1;
  ram[44358]  = 1;
  ram[44359]  = 1;
  ram[44360]  = 1;
  ram[44361]  = 1;
  ram[44362]  = 1;
  ram[44363]  = 1;
  ram[44364]  = 1;
  ram[44365]  = 1;
  ram[44366]  = 1;
  ram[44367]  = 1;
  ram[44368]  = 1;
  ram[44369]  = 1;
  ram[44370]  = 1;
  ram[44371]  = 1;
  ram[44372]  = 1;
  ram[44373]  = 1;
  ram[44374]  = 1;
  ram[44375]  = 1;
  ram[44376]  = 1;
  ram[44377]  = 1;
  ram[44378]  = 1;
  ram[44379]  = 1;
  ram[44380]  = 1;
  ram[44381]  = 1;
  ram[44382]  = 1;
  ram[44383]  = 1;
  ram[44384]  = 1;
  ram[44385]  = 1;
  ram[44386]  = 1;
  ram[44387]  = 1;
  ram[44388]  = 1;
  ram[44389]  = 1;
  ram[44390]  = 1;
  ram[44391]  = 1;
  ram[44392]  = 1;
  ram[44393]  = 1;
  ram[44394]  = 1;
  ram[44395]  = 1;
  ram[44396]  = 1;
  ram[44397]  = 1;
  ram[44398]  = 1;
  ram[44399]  = 1;
  ram[44400]  = 1;
  ram[44401]  = 1;
  ram[44402]  = 1;
  ram[44403]  = 1;
  ram[44404]  = 1;
  ram[44405]  = 1;
  ram[44406]  = 1;
  ram[44407]  = 1;
  ram[44408]  = 1;
  ram[44409]  = 1;
  ram[44410]  = 1;
  ram[44411]  = 1;
  ram[44412]  = 1;
  ram[44413]  = 1;
  ram[44414]  = 1;
  ram[44415]  = 1;
  ram[44416]  = 1;
  ram[44417]  = 1;
  ram[44418]  = 1;
  ram[44419]  = 1;
  ram[44420]  = 1;
  ram[44421]  = 1;
  ram[44422]  = 1;
  ram[44423]  = 1;
  ram[44424]  = 1;
  ram[44425]  = 1;
  ram[44426]  = 1;
  ram[44427]  = 1;
  ram[44428]  = 1;
  ram[44429]  = 1;
  ram[44430]  = 1;
  ram[44431]  = 1;
  ram[44432]  = 1;
  ram[44433]  = 1;
  ram[44434]  = 1;
  ram[44435]  = 1;
  ram[44436]  = 1;
  ram[44437]  = 1;
  ram[44438]  = 1;
  ram[44439]  = 1;
  ram[44440]  = 1;
  ram[44441]  = 1;
  ram[44442]  = 1;
  ram[44443]  = 1;
  ram[44444]  = 1;
  ram[44445]  = 1;
  ram[44446]  = 1;
  ram[44447]  = 1;
  ram[44448]  = 1;
  ram[44449]  = 1;
  ram[44450]  = 1;
  ram[44451]  = 1;
  ram[44452]  = 1;
  ram[44453]  = 1;
  ram[44454]  = 1;
  ram[44455]  = 1;
  ram[44456]  = 1;
  ram[44457]  = 1;
  ram[44458]  = 1;
  ram[44459]  = 1;
  ram[44460]  = 1;
  ram[44461]  = 1;
  ram[44462]  = 1;
  ram[44463]  = 1;
  ram[44464]  = 1;
  ram[44465]  = 1;
  ram[44466]  = 1;
  ram[44467]  = 1;
  ram[44468]  = 1;
  ram[44469]  = 1;
  ram[44470]  = 1;
  ram[44471]  = 1;
  ram[44472]  = 1;
  ram[44473]  = 1;
  ram[44474]  = 1;
  ram[44475]  = 1;
  ram[44476]  = 1;
  ram[44477]  = 1;
  ram[44478]  = 1;
  ram[44479]  = 1;
  ram[44480]  = 1;
  ram[44481]  = 1;
  ram[44482]  = 1;
  ram[44483]  = 1;
  ram[44484]  = 1;
  ram[44485]  = 1;
  ram[44486]  = 1;
  ram[44487]  = 1;
  ram[44488]  = 1;
  ram[44489]  = 1;
  ram[44490]  = 1;
  ram[44491]  = 1;
  ram[44492]  = 1;
  ram[44493]  = 1;
  ram[44494]  = 1;
  ram[44495]  = 1;
  ram[44496]  = 1;
  ram[44497]  = 1;
  ram[44498]  = 1;
  ram[44499]  = 1;
  ram[44500]  = 1;
  ram[44501]  = 1;
  ram[44502]  = 1;
  ram[44503]  = 1;
  ram[44504]  = 1;
  ram[44505]  = 1;
  ram[44506]  = 1;
  ram[44507]  = 1;
  ram[44508]  = 1;
  ram[44509]  = 1;
  ram[44510]  = 1;
  ram[44511]  = 1;
  ram[44512]  = 1;
  ram[44513]  = 1;
  ram[44514]  = 1;
  ram[44515]  = 1;
  ram[44516]  = 1;
  ram[44517]  = 1;
  ram[44518]  = 1;
  ram[44519]  = 1;
  ram[44520]  = 1;
  ram[44521]  = 1;
  ram[44522]  = 1;
  ram[44523]  = 1;
  ram[44524]  = 1;
  ram[44525]  = 1;
  ram[44526]  = 1;
  ram[44527]  = 1;
  ram[44528]  = 1;
  ram[44529]  = 1;
  ram[44530]  = 1;
  ram[44531]  = 1;
  ram[44532]  = 1;
  ram[44533]  = 1;
  ram[44534]  = 1;
  ram[44535]  = 1;
  ram[44536]  = 1;
  ram[44537]  = 1;
  ram[44538]  = 1;
  ram[44539]  = 1;
  ram[44540]  = 1;
  ram[44541]  = 1;
  ram[44542]  = 1;
  ram[44543]  = 1;
  ram[44544]  = 1;
  ram[44545]  = 1;
  ram[44546]  = 1;
  ram[44547]  = 1;
  ram[44548]  = 1;
  ram[44549]  = 1;
  ram[44550]  = 1;
  ram[44551]  = 1;
  ram[44552]  = 1;
  ram[44553]  = 1;
  ram[44554]  = 1;
  ram[44555]  = 1;
  ram[44556]  = 1;
  ram[44557]  = 1;
  ram[44558]  = 1;
  ram[44559]  = 1;
  ram[44560]  = 1;
  ram[44561]  = 1;
  ram[44562]  = 1;
  ram[44563]  = 1;
  ram[44564]  = 1;
  ram[44565]  = 1;
  ram[44566]  = 1;
  ram[44567]  = 1;
  ram[44568]  = 1;
  ram[44569]  = 1;
  ram[44570]  = 1;
  ram[44571]  = 1;
  ram[44572]  = 1;
  ram[44573]  = 1;
  ram[44574]  = 1;
  ram[44575]  = 1;
  ram[44576]  = 1;
  ram[44577]  = 1;
  ram[44578]  = 1;
  ram[44579]  = 1;
  ram[44580]  = 1;
  ram[44581]  = 1;
  ram[44582]  = 1;
  ram[44583]  = 1;
  ram[44584]  = 1;
  ram[44585]  = 1;
  ram[44586]  = 1;
  ram[44587]  = 1;
  ram[44588]  = 1;
  ram[44589]  = 1;
  ram[44590]  = 1;
  ram[44591]  = 1;
  ram[44592]  = 1;
  ram[44593]  = 1;
  ram[44594]  = 1;
  ram[44595]  = 1;
  ram[44596]  = 1;
  ram[44597]  = 1;
  ram[44598]  = 1;
  ram[44599]  = 1;
  ram[44600]  = 1;
  ram[44601]  = 1;
  ram[44602]  = 1;
  ram[44603]  = 1;
  ram[44604]  = 1;
  ram[44605]  = 1;
  ram[44606]  = 1;
  ram[44607]  = 1;
  ram[44608]  = 1;
  ram[44609]  = 1;
  ram[44610]  = 1;
  ram[44611]  = 1;
  ram[44612]  = 1;
  ram[44613]  = 1;
  ram[44614]  = 1;
  ram[44615]  = 1;
  ram[44616]  = 1;
  ram[44617]  = 1;
  ram[44618]  = 1;
  ram[44619]  = 1;
  ram[44620]  = 1;
  ram[44621]  = 1;
  ram[44622]  = 1;
  ram[44623]  = 1;
  ram[44624]  = 1;
  ram[44625]  = 1;
  ram[44626]  = 1;
  ram[44627]  = 1;
  ram[44628]  = 1;
  ram[44629]  = 1;
  ram[44630]  = 1;
  ram[44631]  = 1;
  ram[44632]  = 1;
  ram[44633]  = 1;
  ram[44634]  = 1;
  ram[44635]  = 1;
  ram[44636]  = 1;
  ram[44637]  = 1;
  ram[44638]  = 1;
  ram[44639]  = 1;
  ram[44640]  = 1;
  ram[44641]  = 1;
  ram[44642]  = 1;
  ram[44643]  = 1;
  ram[44644]  = 1;
  ram[44645]  = 1;
  ram[44646]  = 1;
  ram[44647]  = 1;
  ram[44648]  = 1;
  ram[44649]  = 1;
  ram[44650]  = 1;
  ram[44651]  = 1;
  ram[44652]  = 1;
  ram[44653]  = 1;
  ram[44654]  = 1;
  ram[44655]  = 1;
  ram[44656]  = 1;
  ram[44657]  = 1;
  ram[44658]  = 1;
  ram[44659]  = 1;
  ram[44660]  = 1;
  ram[44661]  = 1;
  ram[44662]  = 1;
  ram[44663]  = 1;
  ram[44664]  = 1;
  ram[44665]  = 1;
  ram[44666]  = 1;
  ram[44667]  = 1;
  ram[44668]  = 1;
  ram[44669]  = 1;
  ram[44670]  = 1;
  ram[44671]  = 1;
  ram[44672]  = 1;
  ram[44673]  = 1;
  ram[44674]  = 1;
  ram[44675]  = 1;
  ram[44676]  = 1;
  ram[44677]  = 1;
  ram[44678]  = 1;
  ram[44679]  = 1;
  ram[44680]  = 1;
  ram[44681]  = 1;
  ram[44682]  = 1;
  ram[44683]  = 1;
  ram[44684]  = 1;
  ram[44685]  = 1;
  ram[44686]  = 1;
  ram[44687]  = 1;
  ram[44688]  = 1;
  ram[44689]  = 1;
  ram[44690]  = 1;
  ram[44691]  = 1;
  ram[44692]  = 1;
  ram[44693]  = 1;
  ram[44694]  = 1;
  ram[44695]  = 1;
  ram[44696]  = 1;
  ram[44697]  = 1;
  ram[44698]  = 1;
  ram[44699]  = 1;
  ram[44700]  = 1;
  ram[44701]  = 1;
  ram[44702]  = 1;
  ram[44703]  = 1;
  ram[44704]  = 1;
  ram[44705]  = 1;
  ram[44706]  = 1;
  ram[44707]  = 1;
  ram[44708]  = 1;
  ram[44709]  = 1;
  ram[44710]  = 1;
  ram[44711]  = 1;
  ram[44712]  = 1;
  ram[44713]  = 1;
  ram[44714]  = 1;
  ram[44715]  = 1;
  ram[44716]  = 1;
  ram[44717]  = 1;
  ram[44718]  = 1;
  ram[44719]  = 1;
  ram[44720]  = 1;
  ram[44721]  = 1;
  ram[44722]  = 1;
  ram[44723]  = 1;
  ram[44724]  = 1;
  ram[44725]  = 1;
  ram[44726]  = 1;
  ram[44727]  = 1;
  ram[44728]  = 1;
  ram[44729]  = 1;
  ram[44730]  = 1;
  ram[44731]  = 1;
  ram[44732]  = 1;
  ram[44733]  = 1;
  ram[44734]  = 1;
  ram[44735]  = 1;
  ram[44736]  = 1;
  ram[44737]  = 1;
  ram[44738]  = 1;
  ram[44739]  = 1;
  ram[44740]  = 1;
  ram[44741]  = 1;
  ram[44742]  = 1;
  ram[44743]  = 1;
  ram[44744]  = 1;
  ram[44745]  = 1;
  ram[44746]  = 1;
  ram[44747]  = 1;
  ram[44748]  = 1;
  ram[44749]  = 1;
  ram[44750]  = 1;
  ram[44751]  = 1;
  ram[44752]  = 1;
  ram[44753]  = 1;
  ram[44754]  = 1;
  ram[44755]  = 1;
  ram[44756]  = 1;
  ram[44757]  = 1;
  ram[44758]  = 1;
  ram[44759]  = 1;
  ram[44760]  = 1;
  ram[44761]  = 1;
  ram[44762]  = 1;
  ram[44763]  = 1;
  ram[44764]  = 1;
  ram[44765]  = 1;
  ram[44766]  = 1;
  ram[44767]  = 1;
  ram[44768]  = 1;
  ram[44769]  = 1;
  ram[44770]  = 1;
  ram[44771]  = 1;
  ram[44772]  = 1;
  ram[44773]  = 1;
  ram[44774]  = 1;
  ram[44775]  = 1;
  ram[44776]  = 1;
  ram[44777]  = 1;
  ram[44778]  = 1;
  ram[44779]  = 1;
  ram[44780]  = 1;
  ram[44781]  = 1;
  ram[44782]  = 1;
  ram[44783]  = 1;
  ram[44784]  = 1;
  ram[44785]  = 1;
  ram[44786]  = 1;
  ram[44787]  = 1;
  ram[44788]  = 1;
  ram[44789]  = 1;
  ram[44790]  = 1;
  ram[44791]  = 1;
  ram[44792]  = 1;
  ram[44793]  = 1;
  ram[44794]  = 1;
  ram[44795]  = 1;
  ram[44796]  = 1;
  ram[44797]  = 1;
  ram[44798]  = 1;
  ram[44799]  = 1;
  ram[44800]  = 1;
  ram[44801]  = 1;
  ram[44802]  = 1;
  ram[44803]  = 1;
  ram[44804]  = 1;
  ram[44805]  = 1;
  ram[44806]  = 1;
  ram[44807]  = 1;
  ram[44808]  = 1;
  ram[44809]  = 1;
  ram[44810]  = 1;
  ram[44811]  = 1;
  ram[44812]  = 1;
  ram[44813]  = 1;
  ram[44814]  = 1;
  ram[44815]  = 1;
  ram[44816]  = 1;
  ram[44817]  = 1;
  ram[44818]  = 1;
  ram[44819]  = 1;
  ram[44820]  = 1;
  ram[44821]  = 1;
  ram[44822]  = 1;
  ram[44823]  = 1;
  ram[44824]  = 1;
  ram[44825]  = 1;
  ram[44826]  = 1;
  ram[44827]  = 1;
  ram[44828]  = 1;
  ram[44829]  = 1;
  ram[44830]  = 1;
  ram[44831]  = 1;
  ram[44832]  = 1;
  ram[44833]  = 1;
  ram[44834]  = 1;
  ram[44835]  = 1;
  ram[44836]  = 1;
  ram[44837]  = 1;
  ram[44838]  = 1;
  ram[44839]  = 1;
  ram[44840]  = 1;
  ram[44841]  = 1;
  ram[44842]  = 1;
  ram[44843]  = 1;
  ram[44844]  = 1;
  ram[44845]  = 1;
  ram[44846]  = 1;
  ram[44847]  = 1;
  ram[44848]  = 1;
  ram[44849]  = 1;
  ram[44850]  = 1;
  ram[44851]  = 1;
  ram[44852]  = 1;
  ram[44853]  = 1;
  ram[44854]  = 1;
  ram[44855]  = 1;
  ram[44856]  = 1;
  ram[44857]  = 1;
  ram[44858]  = 1;
  ram[44859]  = 1;
  ram[44860]  = 1;
  ram[44861]  = 1;
  ram[44862]  = 1;
  ram[44863]  = 1;
  ram[44864]  = 1;
  ram[44865]  = 1;
  ram[44866]  = 1;
  ram[44867]  = 1;
  ram[44868]  = 1;
  ram[44869]  = 1;
  ram[44870]  = 1;
  ram[44871]  = 1;
  ram[44872]  = 1;
  ram[44873]  = 1;
  ram[44874]  = 1;
  ram[44875]  = 1;
  ram[44876]  = 1;
  ram[44877]  = 1;
  ram[44878]  = 1;
  ram[44879]  = 1;
  ram[44880]  = 1;
  ram[44881]  = 1;
  ram[44882]  = 1;
  ram[44883]  = 1;
  ram[44884]  = 1;
  ram[44885]  = 1;
  ram[44886]  = 1;
  ram[44887]  = 1;
  ram[44888]  = 1;
  ram[44889]  = 1;
  ram[44890]  = 1;
  ram[44891]  = 1;
  ram[44892]  = 1;
  ram[44893]  = 1;
  ram[44894]  = 1;
  ram[44895]  = 1;
  ram[44896]  = 1;
  ram[44897]  = 1;
  ram[44898]  = 1;
  ram[44899]  = 1;
  ram[44900]  = 1;
  ram[44901]  = 1;
  ram[44902]  = 1;
  ram[44903]  = 1;
  ram[44904]  = 1;
  ram[44905]  = 1;
  ram[44906]  = 1;
  ram[44907]  = 1;
  ram[44908]  = 1;
  ram[44909]  = 1;
  ram[44910]  = 1;
  ram[44911]  = 1;
  ram[44912]  = 1;
  ram[44913]  = 1;
  ram[44914]  = 1;
  ram[44915]  = 1;
  ram[44916]  = 1;
  ram[44917]  = 1;
  ram[44918]  = 1;
  ram[44919]  = 1;
  ram[44920]  = 1;
  ram[44921]  = 1;
  ram[44922]  = 1;
  ram[44923]  = 1;
  ram[44924]  = 1;
  ram[44925]  = 1;
  ram[44926]  = 1;
  ram[44927]  = 1;
  ram[44928]  = 1;
  ram[44929]  = 1;
  ram[44930]  = 1;
  ram[44931]  = 1;
  ram[44932]  = 1;
  ram[44933]  = 1;
  ram[44934]  = 1;
  ram[44935]  = 1;
  ram[44936]  = 1;
  ram[44937]  = 1;
  ram[44938]  = 1;
  ram[44939]  = 1;
  ram[44940]  = 1;
  ram[44941]  = 1;
  ram[44942]  = 1;
  ram[44943]  = 1;
  ram[44944]  = 1;
  ram[44945]  = 1;
  ram[44946]  = 1;
  ram[44947]  = 1;
  ram[44948]  = 1;
  ram[44949]  = 1;
  ram[44950]  = 1;
  ram[44951]  = 1;
  ram[44952]  = 1;
  ram[44953]  = 1;
  ram[44954]  = 1;
  ram[44955]  = 1;
  ram[44956]  = 1;
  ram[44957]  = 1;
  ram[44958]  = 1;
  ram[44959]  = 1;
  ram[44960]  = 1;
  ram[44961]  = 1;
  ram[44962]  = 1;
  ram[44963]  = 1;
  ram[44964]  = 1;
  ram[44965]  = 1;
  ram[44966]  = 1;
  ram[44967]  = 1;
  ram[44968]  = 1;
  ram[44969]  = 1;
  ram[44970]  = 1;
  ram[44971]  = 1;
  ram[44972]  = 1;
  ram[44973]  = 1;
  ram[44974]  = 1;
  ram[44975]  = 1;
  ram[44976]  = 1;
  ram[44977]  = 1;
  ram[44978]  = 1;
  ram[44979]  = 1;
  ram[44980]  = 1;
  ram[44981]  = 1;
  ram[44982]  = 1;
  ram[44983]  = 1;
  ram[44984]  = 1;
  ram[44985]  = 1;
  ram[44986]  = 1;
  ram[44987]  = 1;
  ram[44988]  = 1;
  ram[44989]  = 1;
  ram[44990]  = 1;
  ram[44991]  = 1;
  ram[44992]  = 1;
  ram[44993]  = 1;
  ram[44994]  = 1;
  ram[44995]  = 1;
  ram[44996]  = 1;
  ram[44997]  = 1;
  ram[44998]  = 1;
  ram[44999]  = 1;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
