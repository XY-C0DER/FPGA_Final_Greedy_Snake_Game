module rom_s2 (clock, address, q);
input clock;
output [7:0] q;
input [13:0] address;
reg [7:0] dout;
reg [7:0] ram [16383:0];
assign q = dout;

initial begin
  ram[0]  = 250;
  ram[1]  = 255;
  ram[2]  = 252;
  ram[3]  = 252;
  ram[4]  = 250;
  ram[5]  = 247;
  ram[6]  = 247;
  ram[7]  = 254;
  ram[8]  = 254;
  ram[9]  = 254;
  ram[10]  = 254;
  ram[11]  = 254;
  ram[12]  = 254;
  ram[13]  = 254;
  ram[14]  = 254;
  ram[15]  = 254;
  ram[16]  = 254;
  ram[17]  = 254;
  ram[18]  = 254;
  ram[19]  = 254;
  ram[20]  = 254;
  ram[21]  = 254;
  ram[22]  = 255;
  ram[23]  = 255;
  ram[24]  = 255;
  ram[25]  = 255;
  ram[26]  = 255;
  ram[27]  = 255;
  ram[28]  = 255;
  ram[29]  = 255;
  ram[30]  = 255;
  ram[31]  = 255;
  ram[32]  = 255;
  ram[33]  = 255;
  ram[34]  = 255;
  ram[35]  = 255;
  ram[36]  = 255;
  ram[37]  = 255;
  ram[38]  = 255;
  ram[39]  = 255;
  ram[40]  = 255;
  ram[41]  = 255;
  ram[42]  = 255;
  ram[43]  = 255;
  ram[44]  = 255;
  ram[45]  = 255;
  ram[46]  = 255;
  ram[47]  = 255;
  ram[48]  = 255;
  ram[49]  = 255;
  ram[50]  = 255;
  ram[51]  = 255;
  ram[52]  = 255;
  ram[53]  = 255;
  ram[54]  = 255;
  ram[55]  = 255;
  ram[56]  = 255;
  ram[57]  = 255;
  ram[58]  = 255;
  ram[59]  = 255;
  ram[60]  = 255;
  ram[61]  = 255;
  ram[62]  = 255;
  ram[63]  = 255;
  ram[64]  = 255;
  ram[65]  = 255;
  ram[66]  = 255;
  ram[67]  = 255;
  ram[68]  = 255;
  ram[69]  = 255;
  ram[70]  = 255;
  ram[71]  = 255;
  ram[72]  = 255;
  ram[73]  = 255;
  ram[74]  = 255;
  ram[75]  = 255;
  ram[76]  = 255;
  ram[77]  = 255;
  ram[78]  = 255;
  ram[79]  = 255;
  ram[80]  = 255;
  ram[81]  = 255;
  ram[82]  = 255;
  ram[83]  = 255;
  ram[84]  = 255;
  ram[85]  = 255;
  ram[86]  = 255;
  ram[87]  = 255;
  ram[88]  = 255;
  ram[89]  = 255;
  ram[90]  = 255;
  ram[91]  = 255;
  ram[92]  = 255;
  ram[93]  = 255;
  ram[94]  = 255;
  ram[95]  = 255;
  ram[96]  = 255;
  ram[97]  = 255;
  ram[98]  = 255;
  ram[99]  = 255;
  ram[100]  = 255;
  ram[101]  = 255;
  ram[102]  = 255;
  ram[103]  = 255;
  ram[104]  = 255;
  ram[105]  = 255;
  ram[106]  = 255;
  ram[107]  = 255;
  ram[108]  = 255;
  ram[109]  = 255;
  ram[110]  = 255;
  ram[111]  = 255;
  ram[112]  = 255;
  ram[113]  = 255;
  ram[114]  = 255;
  ram[115]  = 255;
  ram[116]  = 255;
  ram[117]  = 255;
  ram[118]  = 255;
  ram[119]  = 255;
  ram[120]  = 255;
  ram[121]  = 255;
  ram[122]  = 255;
  ram[123]  = 255;
  ram[124]  = 255;
  ram[125]  = 255;
  ram[126]  = 255;
  ram[127]  = 255;
  ram[128]  = 255;
  ram[129]  = 255;
  ram[130]  = 255;
  ram[131]  = 255;
  ram[132]  = 255;
  ram[133]  = 255;
  ram[134]  = 255;
  ram[135]  = 255;
  ram[136]  = 255;
  ram[137]  = 255;
  ram[138]  = 255;
  ram[139]  = 255;
  ram[140]  = 255;
  ram[141]  = 255;
  ram[142]  = 255;
  ram[143]  = 255;
  ram[144]  = 255;
  ram[145]  = 255;
  ram[146]  = 255;
  ram[147]  = 255;
  ram[148]  = 255;
  ram[149]  = 255;
  ram[150]  = 255;
  ram[151]  = 255;
  ram[152]  = 255;
  ram[153]  = 255;
  ram[154]  = 255;
  ram[155]  = 255;
  ram[156]  = 255;
  ram[157]  = 255;
  ram[158]  = 255;
  ram[159]  = 255;
  ram[160]  = 255;
  ram[161]  = 255;
  ram[162]  = 255;
  ram[163]  = 255;
  ram[164]  = 255;
  ram[165]  = 255;
  ram[166]  = 255;
  ram[167]  = 255;
  ram[168]  = 255;
  ram[169]  = 255;
  ram[170]  = 255;
  ram[171]  = 255;
  ram[172]  = 255;
  ram[173]  = 255;
  ram[174]  = 255;
  ram[175]  = 255;
  ram[176]  = 255;
  ram[177]  = 255;
  ram[178]  = 255;
  ram[179]  = 255;
  ram[180]  = 255;
  ram[181]  = 255;
  ram[182]  = 255;
  ram[183]  = 255;
  ram[184]  = 255;
  ram[185]  = 255;
  ram[186]  = 255;
  ram[187]  = 255;
  ram[188]  = 255;
  ram[189]  = 255;
  ram[190]  = 255;
  ram[191]  = 255;
  ram[192]  = 255;
  ram[193]  = 255;
  ram[194]  = 255;
  ram[195]  = 255;
  ram[196]  = 255;
  ram[197]  = 255;
  ram[198]  = 255;
  ram[199]  = 255;
  ram[200]  = 252;
  ram[201]  = 255;
  ram[202]  = 250;
  ram[203]  = 253;
  ram[204]  = 253;
  ram[205]  = 250;
  ram[206]  = 245;
  ram[207]  = 252;
  ram[208]  = 253;
  ram[209]  = 253;
  ram[210]  = 253;
  ram[211]  = 253;
  ram[212]  = 253;
  ram[213]  = 253;
  ram[214]  = 253;
  ram[215]  = 253;
  ram[216]  = 253;
  ram[217]  = 253;
  ram[218]  = 253;
  ram[219]  = 253;
  ram[220]  = 253;
  ram[221]  = 253;
  ram[222]  = 255;
  ram[223]  = 255;
  ram[224]  = 255;
  ram[225]  = 255;
  ram[226]  = 255;
  ram[227]  = 255;
  ram[228]  = 255;
  ram[229]  = 255;
  ram[230]  = 255;
  ram[231]  = 255;
  ram[232]  = 255;
  ram[233]  = 255;
  ram[234]  = 255;
  ram[235]  = 255;
  ram[236]  = 255;
  ram[237]  = 255;
  ram[238]  = 255;
  ram[239]  = 255;
  ram[240]  = 255;
  ram[241]  = 255;
  ram[242]  = 255;
  ram[243]  = 255;
  ram[244]  = 255;
  ram[245]  = 255;
  ram[246]  = 255;
  ram[247]  = 255;
  ram[248]  = 255;
  ram[249]  = 255;
  ram[250]  = 255;
  ram[251]  = 255;
  ram[252]  = 255;
  ram[253]  = 255;
  ram[254]  = 255;
  ram[255]  = 255;
  ram[256]  = 255;
  ram[257]  = 255;
  ram[258]  = 255;
  ram[259]  = 255;
  ram[260]  = 255;
  ram[261]  = 255;
  ram[262]  = 255;
  ram[263]  = 255;
  ram[264]  = 255;
  ram[265]  = 255;
  ram[266]  = 255;
  ram[267]  = 255;
  ram[268]  = 255;
  ram[269]  = 255;
  ram[270]  = 255;
  ram[271]  = 255;
  ram[272]  = 255;
  ram[273]  = 255;
  ram[274]  = 255;
  ram[275]  = 255;
  ram[276]  = 255;
  ram[277]  = 255;
  ram[278]  = 255;
  ram[279]  = 255;
  ram[280]  = 255;
  ram[281]  = 255;
  ram[282]  = 255;
  ram[283]  = 255;
  ram[284]  = 255;
  ram[285]  = 255;
  ram[286]  = 255;
  ram[287]  = 255;
  ram[288]  = 255;
  ram[289]  = 255;
  ram[290]  = 255;
  ram[291]  = 255;
  ram[292]  = 255;
  ram[293]  = 255;
  ram[294]  = 255;
  ram[295]  = 255;
  ram[296]  = 255;
  ram[297]  = 255;
  ram[298]  = 255;
  ram[299]  = 255;
  ram[300]  = 255;
  ram[301]  = 255;
  ram[302]  = 255;
  ram[303]  = 255;
  ram[304]  = 255;
  ram[305]  = 255;
  ram[306]  = 255;
  ram[307]  = 255;
  ram[308]  = 255;
  ram[309]  = 255;
  ram[310]  = 255;
  ram[311]  = 255;
  ram[312]  = 255;
  ram[313]  = 255;
  ram[314]  = 255;
  ram[315]  = 255;
  ram[316]  = 255;
  ram[317]  = 255;
  ram[318]  = 255;
  ram[319]  = 255;
  ram[320]  = 255;
  ram[321]  = 255;
  ram[322]  = 255;
  ram[323]  = 255;
  ram[324]  = 255;
  ram[325]  = 255;
  ram[326]  = 255;
  ram[327]  = 255;
  ram[328]  = 255;
  ram[329]  = 255;
  ram[330]  = 255;
  ram[331]  = 255;
  ram[332]  = 255;
  ram[333]  = 255;
  ram[334]  = 255;
  ram[335]  = 255;
  ram[336]  = 255;
  ram[337]  = 255;
  ram[338]  = 255;
  ram[339]  = 255;
  ram[340]  = 255;
  ram[341]  = 255;
  ram[342]  = 255;
  ram[343]  = 255;
  ram[344]  = 255;
  ram[345]  = 255;
  ram[346]  = 255;
  ram[347]  = 255;
  ram[348]  = 255;
  ram[349]  = 255;
  ram[350]  = 255;
  ram[351]  = 255;
  ram[352]  = 255;
  ram[353]  = 255;
  ram[354]  = 255;
  ram[355]  = 255;
  ram[356]  = 255;
  ram[357]  = 255;
  ram[358]  = 255;
  ram[359]  = 255;
  ram[360]  = 255;
  ram[361]  = 255;
  ram[362]  = 255;
  ram[363]  = 255;
  ram[364]  = 255;
  ram[365]  = 255;
  ram[366]  = 255;
  ram[367]  = 255;
  ram[368]  = 255;
  ram[369]  = 255;
  ram[370]  = 255;
  ram[371]  = 255;
  ram[372]  = 255;
  ram[373]  = 255;
  ram[374]  = 255;
  ram[375]  = 255;
  ram[376]  = 255;
  ram[377]  = 255;
  ram[378]  = 255;
  ram[379]  = 255;
  ram[380]  = 255;
  ram[381]  = 255;
  ram[382]  = 255;
  ram[383]  = 255;
  ram[384]  = 255;
  ram[385]  = 255;
  ram[386]  = 255;
  ram[387]  = 255;
  ram[388]  = 255;
  ram[389]  = 255;
  ram[390]  = 255;
  ram[391]  = 255;
  ram[392]  = 255;
  ram[393]  = 255;
  ram[394]  = 255;
  ram[395]  = 252;
  ram[396]  = 243;
  ram[397]  = 252;
  ram[398]  = 242;
  ram[399]  = 254;
  ram[400]  = 250;
  ram[401]  = 255;
  ram[402]  = 253;
  ram[403]  = 255;
  ram[404]  = 255;
  ram[405]  = 255;
  ram[406]  = 255;
  ram[407]  = 254;
  ram[408]  = 254;
  ram[409]  = 254;
  ram[410]  = 254;
  ram[411]  = 254;
  ram[412]  = 254;
  ram[413]  = 254;
  ram[414]  = 254;
  ram[415]  = 254;
  ram[416]  = 254;
  ram[417]  = 254;
  ram[418]  = 254;
  ram[419]  = 254;
  ram[420]  = 254;
  ram[421]  = 254;
  ram[422]  = 255;
  ram[423]  = 255;
  ram[424]  = 255;
  ram[425]  = 255;
  ram[426]  = 255;
  ram[427]  = 255;
  ram[428]  = 255;
  ram[429]  = 255;
  ram[430]  = 255;
  ram[431]  = 255;
  ram[432]  = 255;
  ram[433]  = 255;
  ram[434]  = 255;
  ram[435]  = 255;
  ram[436]  = 255;
  ram[437]  = 255;
  ram[438]  = 255;
  ram[439]  = 255;
  ram[440]  = 255;
  ram[441]  = 255;
  ram[442]  = 255;
  ram[443]  = 255;
  ram[444]  = 255;
  ram[445]  = 255;
  ram[446]  = 255;
  ram[447]  = 255;
  ram[448]  = 255;
  ram[449]  = 255;
  ram[450]  = 255;
  ram[451]  = 255;
  ram[452]  = 255;
  ram[453]  = 255;
  ram[454]  = 255;
  ram[455]  = 255;
  ram[456]  = 255;
  ram[457]  = 255;
  ram[458]  = 255;
  ram[459]  = 255;
  ram[460]  = 255;
  ram[461]  = 255;
  ram[462]  = 255;
  ram[463]  = 255;
  ram[464]  = 255;
  ram[465]  = 255;
  ram[466]  = 255;
  ram[467]  = 255;
  ram[468]  = 255;
  ram[469]  = 255;
  ram[470]  = 255;
  ram[471]  = 255;
  ram[472]  = 255;
  ram[473]  = 255;
  ram[474]  = 255;
  ram[475]  = 255;
  ram[476]  = 255;
  ram[477]  = 255;
  ram[478]  = 255;
  ram[479]  = 255;
  ram[480]  = 255;
  ram[481]  = 255;
  ram[482]  = 255;
  ram[483]  = 255;
  ram[484]  = 255;
  ram[485]  = 255;
  ram[486]  = 255;
  ram[487]  = 255;
  ram[488]  = 255;
  ram[489]  = 255;
  ram[490]  = 255;
  ram[491]  = 255;
  ram[492]  = 255;
  ram[493]  = 255;
  ram[494]  = 255;
  ram[495]  = 255;
  ram[496]  = 255;
  ram[497]  = 255;
  ram[498]  = 255;
  ram[499]  = 255;
  ram[500]  = 255;
  ram[501]  = 255;
  ram[502]  = 255;
  ram[503]  = 255;
  ram[504]  = 255;
  ram[505]  = 255;
  ram[506]  = 255;
  ram[507]  = 255;
  ram[508]  = 255;
  ram[509]  = 255;
  ram[510]  = 255;
  ram[511]  = 255;
  ram[512]  = 255;
  ram[513]  = 255;
  ram[514]  = 255;
  ram[515]  = 255;
  ram[516]  = 255;
  ram[517]  = 255;
  ram[518]  = 255;
  ram[519]  = 255;
  ram[520]  = 255;
  ram[521]  = 255;
  ram[522]  = 255;
  ram[523]  = 255;
  ram[524]  = 255;
  ram[525]  = 255;
  ram[526]  = 255;
  ram[527]  = 255;
  ram[528]  = 255;
  ram[529]  = 255;
  ram[530]  = 255;
  ram[531]  = 255;
  ram[532]  = 255;
  ram[533]  = 255;
  ram[534]  = 255;
  ram[535]  = 255;
  ram[536]  = 255;
  ram[537]  = 255;
  ram[538]  = 255;
  ram[539]  = 255;
  ram[540]  = 255;
  ram[541]  = 255;
  ram[542]  = 255;
  ram[543]  = 255;
  ram[544]  = 255;
  ram[545]  = 255;
  ram[546]  = 255;
  ram[547]  = 255;
  ram[548]  = 255;
  ram[549]  = 255;
  ram[550]  = 255;
  ram[551]  = 255;
  ram[552]  = 255;
  ram[553]  = 255;
  ram[554]  = 255;
  ram[555]  = 255;
  ram[556]  = 255;
  ram[557]  = 255;
  ram[558]  = 255;
  ram[559]  = 255;
  ram[560]  = 255;
  ram[561]  = 255;
  ram[562]  = 255;
  ram[563]  = 255;
  ram[564]  = 255;
  ram[565]  = 255;
  ram[566]  = 255;
  ram[567]  = 255;
  ram[568]  = 255;
  ram[569]  = 255;
  ram[570]  = 255;
  ram[571]  = 255;
  ram[572]  = 255;
  ram[573]  = 255;
  ram[574]  = 255;
  ram[575]  = 255;
  ram[576]  = 255;
  ram[577]  = 255;
  ram[578]  = 255;
  ram[579]  = 255;
  ram[580]  = 255;
  ram[581]  = 255;
  ram[582]  = 255;
  ram[583]  = 255;
  ram[584]  = 255;
  ram[585]  = 255;
  ram[586]  = 255;
  ram[587]  = 255;
  ram[588]  = 255;
  ram[589]  = 255;
  ram[590]  = 255;
  ram[591]  = 255;
  ram[592]  = 255;
  ram[593]  = 255;
  ram[594]  = 255;
  ram[595]  = 255;
  ram[596]  = 252;
  ram[597]  = 255;
  ram[598]  = 242;
  ram[599]  = 254;
  ram[600]  = 254;
  ram[601]  = 228;
  ram[602]  = 199;
  ram[603]  = 219;
  ram[604]  = 217;
  ram[605]  = 222;
  ram[606]  = 227;
  ram[607]  = 224;
  ram[608]  = 224;
  ram[609]  = 224;
  ram[610]  = 224;
  ram[611]  = 224;
  ram[612]  = 224;
  ram[613]  = 224;
  ram[614]  = 224;
  ram[615]  = 224;
  ram[616]  = 224;
  ram[617]  = 224;
  ram[618]  = 224;
  ram[619]  = 224;
  ram[620]  = 224;
  ram[621]  = 224;
  ram[622]  = 223;
  ram[623]  = 223;
  ram[624]  = 223;
  ram[625]  = 223;
  ram[626]  = 223;
  ram[627]  = 223;
  ram[628]  = 223;
  ram[629]  = 223;
  ram[630]  = 223;
  ram[631]  = 223;
  ram[632]  = 223;
  ram[633]  = 223;
  ram[634]  = 223;
  ram[635]  = 223;
  ram[636]  = 223;
  ram[637]  = 223;
  ram[638]  = 223;
  ram[639]  = 223;
  ram[640]  = 223;
  ram[641]  = 223;
  ram[642]  = 223;
  ram[643]  = 223;
  ram[644]  = 223;
  ram[645]  = 223;
  ram[646]  = 223;
  ram[647]  = 223;
  ram[648]  = 223;
  ram[649]  = 223;
  ram[650]  = 223;
  ram[651]  = 223;
  ram[652]  = 223;
  ram[653]  = 223;
  ram[654]  = 223;
  ram[655]  = 223;
  ram[656]  = 223;
  ram[657]  = 223;
  ram[658]  = 223;
  ram[659]  = 223;
  ram[660]  = 223;
  ram[661]  = 223;
  ram[662]  = 223;
  ram[663]  = 223;
  ram[664]  = 223;
  ram[665]  = 223;
  ram[666]  = 223;
  ram[667]  = 223;
  ram[668]  = 223;
  ram[669]  = 223;
  ram[670]  = 223;
  ram[671]  = 223;
  ram[672]  = 223;
  ram[673]  = 223;
  ram[674]  = 223;
  ram[675]  = 223;
  ram[676]  = 223;
  ram[677]  = 223;
  ram[678]  = 223;
  ram[679]  = 223;
  ram[680]  = 223;
  ram[681]  = 223;
  ram[682]  = 223;
  ram[683]  = 223;
  ram[684]  = 223;
  ram[685]  = 223;
  ram[686]  = 223;
  ram[687]  = 223;
  ram[688]  = 223;
  ram[689]  = 223;
  ram[690]  = 223;
  ram[691]  = 223;
  ram[692]  = 223;
  ram[693]  = 223;
  ram[694]  = 223;
  ram[695]  = 223;
  ram[696]  = 223;
  ram[697]  = 223;
  ram[698]  = 223;
  ram[699]  = 223;
  ram[700]  = 223;
  ram[701]  = 223;
  ram[702]  = 223;
  ram[703]  = 223;
  ram[704]  = 223;
  ram[705]  = 223;
  ram[706]  = 223;
  ram[707]  = 223;
  ram[708]  = 223;
  ram[709]  = 223;
  ram[710]  = 223;
  ram[711]  = 223;
  ram[712]  = 223;
  ram[713]  = 223;
  ram[714]  = 223;
  ram[715]  = 223;
  ram[716]  = 223;
  ram[717]  = 223;
  ram[718]  = 223;
  ram[719]  = 223;
  ram[720]  = 223;
  ram[721]  = 223;
  ram[722]  = 223;
  ram[723]  = 223;
  ram[724]  = 223;
  ram[725]  = 223;
  ram[726]  = 223;
  ram[727]  = 223;
  ram[728]  = 223;
  ram[729]  = 223;
  ram[730]  = 223;
  ram[731]  = 223;
  ram[732]  = 223;
  ram[733]  = 223;
  ram[734]  = 223;
  ram[735]  = 223;
  ram[736]  = 223;
  ram[737]  = 223;
  ram[738]  = 223;
  ram[739]  = 223;
  ram[740]  = 223;
  ram[741]  = 223;
  ram[742]  = 223;
  ram[743]  = 223;
  ram[744]  = 223;
  ram[745]  = 223;
  ram[746]  = 223;
  ram[747]  = 223;
  ram[748]  = 223;
  ram[749]  = 223;
  ram[750]  = 223;
  ram[751]  = 223;
  ram[752]  = 223;
  ram[753]  = 223;
  ram[754]  = 223;
  ram[755]  = 223;
  ram[756]  = 223;
  ram[757]  = 223;
  ram[758]  = 223;
  ram[759]  = 223;
  ram[760]  = 223;
  ram[761]  = 223;
  ram[762]  = 223;
  ram[763]  = 223;
  ram[764]  = 223;
  ram[765]  = 223;
  ram[766]  = 223;
  ram[767]  = 223;
  ram[768]  = 223;
  ram[769]  = 223;
  ram[770]  = 223;
  ram[771]  = 223;
  ram[772]  = 223;
  ram[773]  = 223;
  ram[774]  = 223;
  ram[775]  = 223;
  ram[776]  = 223;
  ram[777]  = 223;
  ram[778]  = 223;
  ram[779]  = 223;
  ram[780]  = 223;
  ram[781]  = 223;
  ram[782]  = 223;
  ram[783]  = 223;
  ram[784]  = 223;
  ram[785]  = 223;
  ram[786]  = 223;
  ram[787]  = 223;
  ram[788]  = 223;
  ram[789]  = 223;
  ram[790]  = 223;
  ram[791]  = 223;
  ram[792]  = 223;
  ram[793]  = 223;
  ram[794]  = 223;
  ram[795]  = 220;
  ram[796]  = 210;
  ram[797]  = 206;
  ram[798]  = 245;
  ram[799]  = 255;
  ram[800]  = 254;
  ram[801]  = 230;
  ram[802]  = 219;
  ram[803]  = 221;
  ram[804]  = 201;
  ram[805]  = 200;
  ram[806]  = 209;
  ram[807]  = 209;
  ram[808]  = 209;
  ram[809]  = 209;
  ram[810]  = 209;
  ram[811]  = 209;
  ram[812]  = 209;
  ram[813]  = 209;
  ram[814]  = 209;
  ram[815]  = 209;
  ram[816]  = 209;
  ram[817]  = 209;
  ram[818]  = 209;
  ram[819]  = 209;
  ram[820]  = 209;
  ram[821]  = 208;
  ram[822]  = 203;
  ram[823]  = 203;
  ram[824]  = 203;
  ram[825]  = 203;
  ram[826]  = 203;
  ram[827]  = 203;
  ram[828]  = 203;
  ram[829]  = 203;
  ram[830]  = 203;
  ram[831]  = 203;
  ram[832]  = 203;
  ram[833]  = 203;
  ram[834]  = 203;
  ram[835]  = 203;
  ram[836]  = 203;
  ram[837]  = 203;
  ram[838]  = 203;
  ram[839]  = 203;
  ram[840]  = 203;
  ram[841]  = 203;
  ram[842]  = 203;
  ram[843]  = 203;
  ram[844]  = 203;
  ram[845]  = 203;
  ram[846]  = 203;
  ram[847]  = 203;
  ram[848]  = 203;
  ram[849]  = 203;
  ram[850]  = 203;
  ram[851]  = 203;
  ram[852]  = 203;
  ram[853]  = 203;
  ram[854]  = 203;
  ram[855]  = 203;
  ram[856]  = 203;
  ram[857]  = 203;
  ram[858]  = 203;
  ram[859]  = 203;
  ram[860]  = 203;
  ram[861]  = 203;
  ram[862]  = 203;
  ram[863]  = 203;
  ram[864]  = 203;
  ram[865]  = 203;
  ram[866]  = 203;
  ram[867]  = 203;
  ram[868]  = 203;
  ram[869]  = 203;
  ram[870]  = 203;
  ram[871]  = 203;
  ram[872]  = 203;
  ram[873]  = 203;
  ram[874]  = 203;
  ram[875]  = 203;
  ram[876]  = 203;
  ram[877]  = 203;
  ram[878]  = 203;
  ram[879]  = 203;
  ram[880]  = 203;
  ram[881]  = 203;
  ram[882]  = 203;
  ram[883]  = 203;
  ram[884]  = 203;
  ram[885]  = 203;
  ram[886]  = 203;
  ram[887]  = 203;
  ram[888]  = 203;
  ram[889]  = 203;
  ram[890]  = 203;
  ram[891]  = 203;
  ram[892]  = 203;
  ram[893]  = 203;
  ram[894]  = 203;
  ram[895]  = 203;
  ram[896]  = 203;
  ram[897]  = 203;
  ram[898]  = 203;
  ram[899]  = 203;
  ram[900]  = 203;
  ram[901]  = 203;
  ram[902]  = 203;
  ram[903]  = 203;
  ram[904]  = 203;
  ram[905]  = 203;
  ram[906]  = 203;
  ram[907]  = 203;
  ram[908]  = 203;
  ram[909]  = 203;
  ram[910]  = 203;
  ram[911]  = 203;
  ram[912]  = 203;
  ram[913]  = 203;
  ram[914]  = 203;
  ram[915]  = 203;
  ram[916]  = 203;
  ram[917]  = 203;
  ram[918]  = 203;
  ram[919]  = 203;
  ram[920]  = 203;
  ram[921]  = 203;
  ram[922]  = 203;
  ram[923]  = 203;
  ram[924]  = 203;
  ram[925]  = 203;
  ram[926]  = 203;
  ram[927]  = 203;
  ram[928]  = 203;
  ram[929]  = 203;
  ram[930]  = 203;
  ram[931]  = 203;
  ram[932]  = 203;
  ram[933]  = 203;
  ram[934]  = 203;
  ram[935]  = 203;
  ram[936]  = 203;
  ram[937]  = 203;
  ram[938]  = 203;
  ram[939]  = 203;
  ram[940]  = 203;
  ram[941]  = 203;
  ram[942]  = 203;
  ram[943]  = 203;
  ram[944]  = 203;
  ram[945]  = 203;
  ram[946]  = 203;
  ram[947]  = 203;
  ram[948]  = 203;
  ram[949]  = 203;
  ram[950]  = 203;
  ram[951]  = 203;
  ram[952]  = 203;
  ram[953]  = 203;
  ram[954]  = 203;
  ram[955]  = 203;
  ram[956]  = 203;
  ram[957]  = 203;
  ram[958]  = 203;
  ram[959]  = 203;
  ram[960]  = 203;
  ram[961]  = 203;
  ram[962]  = 203;
  ram[963]  = 203;
  ram[964]  = 203;
  ram[965]  = 203;
  ram[966]  = 203;
  ram[967]  = 203;
  ram[968]  = 203;
  ram[969]  = 203;
  ram[970]  = 203;
  ram[971]  = 203;
  ram[972]  = 203;
  ram[973]  = 203;
  ram[974]  = 203;
  ram[975]  = 203;
  ram[976]  = 203;
  ram[977]  = 203;
  ram[978]  = 203;
  ram[979]  = 203;
  ram[980]  = 203;
  ram[981]  = 203;
  ram[982]  = 203;
  ram[983]  = 203;
  ram[984]  = 203;
  ram[985]  = 203;
  ram[986]  = 203;
  ram[987]  = 203;
  ram[988]  = 203;
  ram[989]  = 203;
  ram[990]  = 203;
  ram[991]  = 203;
  ram[992]  = 203;
  ram[993]  = 203;
  ram[994]  = 203;
  ram[995]  = 201;
  ram[996]  = 219;
  ram[997]  = 216;
  ram[998]  = 244;
  ram[999]  = 255;
  ram[1000]  = 255;
  ram[1001]  = 233;
  ram[1002]  = 201;
  ram[1003]  = 235;
  ram[1004]  = 243;
  ram[1005]  = 241;
  ram[1006]  = 242;
  ram[1007]  = 241;
  ram[1008]  = 241;
  ram[1009]  = 241;
  ram[1010]  = 241;
  ram[1011]  = 241;
  ram[1012]  = 241;
  ram[1013]  = 241;
  ram[1014]  = 241;
  ram[1015]  = 241;
  ram[1016]  = 241;
  ram[1017]  = 241;
  ram[1018]  = 241;
  ram[1019]  = 241;
  ram[1020]  = 242;
  ram[1021]  = 241;
  ram[1022]  = 241;
  ram[1023]  = 241;
  ram[1024]  = 241;
  ram[1025]  = 241;
  ram[1026]  = 241;
  ram[1027]  = 241;
  ram[1028]  = 241;
  ram[1029]  = 241;
  ram[1030]  = 241;
  ram[1031]  = 241;
  ram[1032]  = 241;
  ram[1033]  = 241;
  ram[1034]  = 241;
  ram[1035]  = 241;
  ram[1036]  = 241;
  ram[1037]  = 241;
  ram[1038]  = 241;
  ram[1039]  = 241;
  ram[1040]  = 241;
  ram[1041]  = 241;
  ram[1042]  = 241;
  ram[1043]  = 241;
  ram[1044]  = 241;
  ram[1045]  = 241;
  ram[1046]  = 241;
  ram[1047]  = 241;
  ram[1048]  = 241;
  ram[1049]  = 241;
  ram[1050]  = 241;
  ram[1051]  = 241;
  ram[1052]  = 241;
  ram[1053]  = 241;
  ram[1054]  = 241;
  ram[1055]  = 241;
  ram[1056]  = 241;
  ram[1057]  = 241;
  ram[1058]  = 241;
  ram[1059]  = 241;
  ram[1060]  = 241;
  ram[1061]  = 241;
  ram[1062]  = 241;
  ram[1063]  = 241;
  ram[1064]  = 241;
  ram[1065]  = 241;
  ram[1066]  = 241;
  ram[1067]  = 241;
  ram[1068]  = 241;
  ram[1069]  = 241;
  ram[1070]  = 241;
  ram[1071]  = 241;
  ram[1072]  = 241;
  ram[1073]  = 241;
  ram[1074]  = 241;
  ram[1075]  = 241;
  ram[1076]  = 241;
  ram[1077]  = 241;
  ram[1078]  = 241;
  ram[1079]  = 241;
  ram[1080]  = 241;
  ram[1081]  = 241;
  ram[1082]  = 241;
  ram[1083]  = 241;
  ram[1084]  = 241;
  ram[1085]  = 241;
  ram[1086]  = 241;
  ram[1087]  = 241;
  ram[1088]  = 241;
  ram[1089]  = 241;
  ram[1090]  = 241;
  ram[1091]  = 241;
  ram[1092]  = 241;
  ram[1093]  = 241;
  ram[1094]  = 241;
  ram[1095]  = 241;
  ram[1096]  = 241;
  ram[1097]  = 241;
  ram[1098]  = 241;
  ram[1099]  = 241;
  ram[1100]  = 241;
  ram[1101]  = 241;
  ram[1102]  = 241;
  ram[1103]  = 241;
  ram[1104]  = 241;
  ram[1105]  = 241;
  ram[1106]  = 241;
  ram[1107]  = 241;
  ram[1108]  = 241;
  ram[1109]  = 241;
  ram[1110]  = 241;
  ram[1111]  = 241;
  ram[1112]  = 241;
  ram[1113]  = 241;
  ram[1114]  = 241;
  ram[1115]  = 241;
  ram[1116]  = 241;
  ram[1117]  = 241;
  ram[1118]  = 241;
  ram[1119]  = 241;
  ram[1120]  = 241;
  ram[1121]  = 241;
  ram[1122]  = 241;
  ram[1123]  = 241;
  ram[1124]  = 241;
  ram[1125]  = 241;
  ram[1126]  = 241;
  ram[1127]  = 241;
  ram[1128]  = 241;
  ram[1129]  = 241;
  ram[1130]  = 241;
  ram[1131]  = 241;
  ram[1132]  = 241;
  ram[1133]  = 241;
  ram[1134]  = 241;
  ram[1135]  = 241;
  ram[1136]  = 241;
  ram[1137]  = 241;
  ram[1138]  = 241;
  ram[1139]  = 241;
  ram[1140]  = 241;
  ram[1141]  = 241;
  ram[1142]  = 241;
  ram[1143]  = 241;
  ram[1144]  = 241;
  ram[1145]  = 241;
  ram[1146]  = 241;
  ram[1147]  = 241;
  ram[1148]  = 241;
  ram[1149]  = 241;
  ram[1150]  = 241;
  ram[1151]  = 241;
  ram[1152]  = 241;
  ram[1153]  = 241;
  ram[1154]  = 241;
  ram[1155]  = 241;
  ram[1156]  = 241;
  ram[1157]  = 241;
  ram[1158]  = 241;
  ram[1159]  = 241;
  ram[1160]  = 241;
  ram[1161]  = 241;
  ram[1162]  = 241;
  ram[1163]  = 241;
  ram[1164]  = 241;
  ram[1165]  = 241;
  ram[1166]  = 241;
  ram[1167]  = 241;
  ram[1168]  = 241;
  ram[1169]  = 241;
  ram[1170]  = 241;
  ram[1171]  = 241;
  ram[1172]  = 241;
  ram[1173]  = 241;
  ram[1174]  = 241;
  ram[1175]  = 241;
  ram[1176]  = 241;
  ram[1177]  = 241;
  ram[1178]  = 241;
  ram[1179]  = 241;
  ram[1180]  = 241;
  ram[1181]  = 241;
  ram[1182]  = 241;
  ram[1183]  = 241;
  ram[1184]  = 241;
  ram[1185]  = 241;
  ram[1186]  = 241;
  ram[1187]  = 241;
  ram[1188]  = 241;
  ram[1189]  = 241;
  ram[1190]  = 241;
  ram[1191]  = 241;
  ram[1192]  = 241;
  ram[1193]  = 241;
  ram[1194]  = 241;
  ram[1195]  = 242;
  ram[1196]  = 231;
  ram[1197]  = 203;
  ram[1198]  = 241;
  ram[1199]  = 255;
  ram[1200]  = 255;
  ram[1201]  = 234;
  ram[1202]  = 208;
  ram[1203]  = 245;
  ram[1204]  = 255;
  ram[1205]  = 255;
  ram[1206]  = 254;
  ram[1207]  = 255;
  ram[1208]  = 255;
  ram[1209]  = 255;
  ram[1210]  = 255;
  ram[1211]  = 255;
  ram[1212]  = 255;
  ram[1213]  = 255;
  ram[1214]  = 255;
  ram[1215]  = 255;
  ram[1216]  = 255;
  ram[1217]  = 255;
  ram[1218]  = 255;
  ram[1219]  = 255;
  ram[1220]  = 255;
  ram[1221]  = 255;
  ram[1222]  = 255;
  ram[1223]  = 255;
  ram[1224]  = 255;
  ram[1225]  = 255;
  ram[1226]  = 255;
  ram[1227]  = 255;
  ram[1228]  = 255;
  ram[1229]  = 255;
  ram[1230]  = 255;
  ram[1231]  = 255;
  ram[1232]  = 255;
  ram[1233]  = 255;
  ram[1234]  = 255;
  ram[1235]  = 255;
  ram[1236]  = 255;
  ram[1237]  = 255;
  ram[1238]  = 255;
  ram[1239]  = 255;
  ram[1240]  = 255;
  ram[1241]  = 255;
  ram[1242]  = 255;
  ram[1243]  = 255;
  ram[1244]  = 255;
  ram[1245]  = 255;
  ram[1246]  = 255;
  ram[1247]  = 255;
  ram[1248]  = 255;
  ram[1249]  = 255;
  ram[1250]  = 255;
  ram[1251]  = 255;
  ram[1252]  = 255;
  ram[1253]  = 255;
  ram[1254]  = 255;
  ram[1255]  = 255;
  ram[1256]  = 255;
  ram[1257]  = 255;
  ram[1258]  = 255;
  ram[1259]  = 255;
  ram[1260]  = 255;
  ram[1261]  = 255;
  ram[1262]  = 255;
  ram[1263]  = 255;
  ram[1264]  = 255;
  ram[1265]  = 255;
  ram[1266]  = 255;
  ram[1267]  = 255;
  ram[1268]  = 255;
  ram[1269]  = 255;
  ram[1270]  = 255;
  ram[1271]  = 255;
  ram[1272]  = 255;
  ram[1273]  = 255;
  ram[1274]  = 255;
  ram[1275]  = 255;
  ram[1276]  = 255;
  ram[1277]  = 255;
  ram[1278]  = 255;
  ram[1279]  = 255;
  ram[1280]  = 255;
  ram[1281]  = 255;
  ram[1282]  = 255;
  ram[1283]  = 255;
  ram[1284]  = 255;
  ram[1285]  = 255;
  ram[1286]  = 255;
  ram[1287]  = 255;
  ram[1288]  = 255;
  ram[1289]  = 255;
  ram[1290]  = 255;
  ram[1291]  = 255;
  ram[1292]  = 255;
  ram[1293]  = 255;
  ram[1294]  = 255;
  ram[1295]  = 255;
  ram[1296]  = 255;
  ram[1297]  = 255;
  ram[1298]  = 255;
  ram[1299]  = 255;
  ram[1300]  = 255;
  ram[1301]  = 255;
  ram[1302]  = 255;
  ram[1303]  = 255;
  ram[1304]  = 255;
  ram[1305]  = 255;
  ram[1306]  = 255;
  ram[1307]  = 255;
  ram[1308]  = 255;
  ram[1309]  = 255;
  ram[1310]  = 255;
  ram[1311]  = 255;
  ram[1312]  = 255;
  ram[1313]  = 255;
  ram[1314]  = 255;
  ram[1315]  = 255;
  ram[1316]  = 255;
  ram[1317]  = 255;
  ram[1318]  = 255;
  ram[1319]  = 255;
  ram[1320]  = 255;
  ram[1321]  = 255;
  ram[1322]  = 255;
  ram[1323]  = 255;
  ram[1324]  = 255;
  ram[1325]  = 255;
  ram[1326]  = 255;
  ram[1327]  = 255;
  ram[1328]  = 255;
  ram[1329]  = 255;
  ram[1330]  = 255;
  ram[1331]  = 255;
  ram[1332]  = 255;
  ram[1333]  = 255;
  ram[1334]  = 255;
  ram[1335]  = 255;
  ram[1336]  = 255;
  ram[1337]  = 255;
  ram[1338]  = 255;
  ram[1339]  = 255;
  ram[1340]  = 255;
  ram[1341]  = 255;
  ram[1342]  = 255;
  ram[1343]  = 255;
  ram[1344]  = 255;
  ram[1345]  = 255;
  ram[1346]  = 255;
  ram[1347]  = 255;
  ram[1348]  = 255;
  ram[1349]  = 255;
  ram[1350]  = 255;
  ram[1351]  = 255;
  ram[1352]  = 255;
  ram[1353]  = 255;
  ram[1354]  = 255;
  ram[1355]  = 255;
  ram[1356]  = 255;
  ram[1357]  = 255;
  ram[1358]  = 255;
  ram[1359]  = 255;
  ram[1360]  = 255;
  ram[1361]  = 255;
  ram[1362]  = 255;
  ram[1363]  = 255;
  ram[1364]  = 255;
  ram[1365]  = 255;
  ram[1366]  = 255;
  ram[1367]  = 255;
  ram[1368]  = 255;
  ram[1369]  = 255;
  ram[1370]  = 255;
  ram[1371]  = 255;
  ram[1372]  = 255;
  ram[1373]  = 255;
  ram[1374]  = 255;
  ram[1375]  = 255;
  ram[1376]  = 255;
  ram[1377]  = 255;
  ram[1378]  = 255;
  ram[1379]  = 255;
  ram[1380]  = 255;
  ram[1381]  = 255;
  ram[1382]  = 255;
  ram[1383]  = 255;
  ram[1384]  = 255;
  ram[1385]  = 255;
  ram[1386]  = 255;
  ram[1387]  = 255;
  ram[1388]  = 255;
  ram[1389]  = 255;
  ram[1390]  = 255;
  ram[1391]  = 255;
  ram[1392]  = 255;
  ram[1393]  = 255;
  ram[1394]  = 255;
  ram[1395]  = 255;
  ram[1396]  = 236;
  ram[1397]  = 212;
  ram[1398]  = 243;
  ram[1399]  = 255;
  ram[1400]  = 255;
  ram[1401]  = 234;
  ram[1402]  = 208;
  ram[1403]  = 244;
  ram[1404]  = 255;
  ram[1405]  = 254;
  ram[1406]  = 252;
  ram[1407]  = 255;
  ram[1408]  = 255;
  ram[1409]  = 255;
  ram[1410]  = 255;
  ram[1411]  = 255;
  ram[1412]  = 255;
  ram[1413]  = 255;
  ram[1414]  = 255;
  ram[1415]  = 255;
  ram[1416]  = 255;
  ram[1417]  = 255;
  ram[1418]  = 255;
  ram[1419]  = 255;
  ram[1420]  = 255;
  ram[1421]  = 255;
  ram[1422]  = 255;
  ram[1423]  = 255;
  ram[1424]  = 255;
  ram[1425]  = 255;
  ram[1426]  = 255;
  ram[1427]  = 255;
  ram[1428]  = 255;
  ram[1429]  = 255;
  ram[1430]  = 255;
  ram[1431]  = 255;
  ram[1432]  = 255;
  ram[1433]  = 255;
  ram[1434]  = 255;
  ram[1435]  = 255;
  ram[1436]  = 255;
  ram[1437]  = 255;
  ram[1438]  = 255;
  ram[1439]  = 255;
  ram[1440]  = 255;
  ram[1441]  = 255;
  ram[1442]  = 255;
  ram[1443]  = 255;
  ram[1444]  = 255;
  ram[1445]  = 255;
  ram[1446]  = 255;
  ram[1447]  = 255;
  ram[1448]  = 255;
  ram[1449]  = 255;
  ram[1450]  = 255;
  ram[1451]  = 255;
  ram[1452]  = 255;
  ram[1453]  = 255;
  ram[1454]  = 255;
  ram[1455]  = 255;
  ram[1456]  = 255;
  ram[1457]  = 255;
  ram[1458]  = 255;
  ram[1459]  = 255;
  ram[1460]  = 255;
  ram[1461]  = 255;
  ram[1462]  = 255;
  ram[1463]  = 255;
  ram[1464]  = 255;
  ram[1465]  = 255;
  ram[1466]  = 255;
  ram[1467]  = 255;
  ram[1468]  = 255;
  ram[1469]  = 255;
  ram[1470]  = 255;
  ram[1471]  = 255;
  ram[1472]  = 255;
  ram[1473]  = 255;
  ram[1474]  = 255;
  ram[1475]  = 255;
  ram[1476]  = 255;
  ram[1477]  = 255;
  ram[1478]  = 255;
  ram[1479]  = 255;
  ram[1480]  = 255;
  ram[1481]  = 255;
  ram[1482]  = 255;
  ram[1483]  = 255;
  ram[1484]  = 255;
  ram[1485]  = 255;
  ram[1486]  = 255;
  ram[1487]  = 255;
  ram[1488]  = 255;
  ram[1489]  = 255;
  ram[1490]  = 255;
  ram[1491]  = 255;
  ram[1492]  = 255;
  ram[1493]  = 255;
  ram[1494]  = 255;
  ram[1495]  = 255;
  ram[1496]  = 255;
  ram[1497]  = 255;
  ram[1498]  = 255;
  ram[1499]  = 255;
  ram[1500]  = 255;
  ram[1501]  = 255;
  ram[1502]  = 255;
  ram[1503]  = 255;
  ram[1504]  = 255;
  ram[1505]  = 255;
  ram[1506]  = 255;
  ram[1507]  = 255;
  ram[1508]  = 255;
  ram[1509]  = 255;
  ram[1510]  = 255;
  ram[1511]  = 255;
  ram[1512]  = 255;
  ram[1513]  = 255;
  ram[1514]  = 255;
  ram[1515]  = 255;
  ram[1516]  = 255;
  ram[1517]  = 255;
  ram[1518]  = 255;
  ram[1519]  = 255;
  ram[1520]  = 255;
  ram[1521]  = 255;
  ram[1522]  = 255;
  ram[1523]  = 255;
  ram[1524]  = 255;
  ram[1525]  = 255;
  ram[1526]  = 255;
  ram[1527]  = 255;
  ram[1528]  = 255;
  ram[1529]  = 255;
  ram[1530]  = 255;
  ram[1531]  = 255;
  ram[1532]  = 255;
  ram[1533]  = 255;
  ram[1534]  = 255;
  ram[1535]  = 255;
  ram[1536]  = 255;
  ram[1537]  = 255;
  ram[1538]  = 255;
  ram[1539]  = 255;
  ram[1540]  = 255;
  ram[1541]  = 255;
  ram[1542]  = 255;
  ram[1543]  = 255;
  ram[1544]  = 255;
  ram[1545]  = 255;
  ram[1546]  = 255;
  ram[1547]  = 255;
  ram[1548]  = 255;
  ram[1549]  = 255;
  ram[1550]  = 255;
  ram[1551]  = 255;
  ram[1552]  = 255;
  ram[1553]  = 255;
  ram[1554]  = 255;
  ram[1555]  = 255;
  ram[1556]  = 255;
  ram[1557]  = 255;
  ram[1558]  = 255;
  ram[1559]  = 255;
  ram[1560]  = 255;
  ram[1561]  = 255;
  ram[1562]  = 255;
  ram[1563]  = 255;
  ram[1564]  = 255;
  ram[1565]  = 255;
  ram[1566]  = 255;
  ram[1567]  = 255;
  ram[1568]  = 255;
  ram[1569]  = 255;
  ram[1570]  = 255;
  ram[1571]  = 255;
  ram[1572]  = 255;
  ram[1573]  = 255;
  ram[1574]  = 255;
  ram[1575]  = 255;
  ram[1576]  = 255;
  ram[1577]  = 255;
  ram[1578]  = 255;
  ram[1579]  = 255;
  ram[1580]  = 255;
  ram[1581]  = 255;
  ram[1582]  = 255;
  ram[1583]  = 255;
  ram[1584]  = 255;
  ram[1585]  = 255;
  ram[1586]  = 255;
  ram[1587]  = 255;
  ram[1588]  = 255;
  ram[1589]  = 255;
  ram[1590]  = 255;
  ram[1591]  = 255;
  ram[1592]  = 255;
  ram[1593]  = 255;
  ram[1594]  = 255;
  ram[1595]  = 255;
  ram[1596]  = 236;
  ram[1597]  = 211;
  ram[1598]  = 243;
  ram[1599]  = 255;
  ram[1600]  = 255;
  ram[1601]  = 234;
  ram[1602]  = 207;
  ram[1603]  = 243;
  ram[1604]  = 255;
  ram[1605]  = 254;
  ram[1606]  = 252;
  ram[1607]  = 255;
  ram[1608]  = 255;
  ram[1609]  = 255;
  ram[1610]  = 255;
  ram[1611]  = 255;
  ram[1612]  = 255;
  ram[1613]  = 255;
  ram[1614]  = 255;
  ram[1615]  = 255;
  ram[1616]  = 255;
  ram[1617]  = 255;
  ram[1618]  = 255;
  ram[1619]  = 255;
  ram[1620]  = 255;
  ram[1621]  = 255;
  ram[1622]  = 255;
  ram[1623]  = 255;
  ram[1624]  = 255;
  ram[1625]  = 255;
  ram[1626]  = 255;
  ram[1627]  = 255;
  ram[1628]  = 255;
  ram[1629]  = 255;
  ram[1630]  = 255;
  ram[1631]  = 255;
  ram[1632]  = 255;
  ram[1633]  = 255;
  ram[1634]  = 255;
  ram[1635]  = 255;
  ram[1636]  = 255;
  ram[1637]  = 255;
  ram[1638]  = 255;
  ram[1639]  = 255;
  ram[1640]  = 255;
  ram[1641]  = 255;
  ram[1642]  = 255;
  ram[1643]  = 255;
  ram[1644]  = 255;
  ram[1645]  = 255;
  ram[1646]  = 255;
  ram[1647]  = 255;
  ram[1648]  = 255;
  ram[1649]  = 255;
  ram[1650]  = 255;
  ram[1651]  = 255;
  ram[1652]  = 255;
  ram[1653]  = 255;
  ram[1654]  = 255;
  ram[1655]  = 255;
  ram[1656]  = 255;
  ram[1657]  = 255;
  ram[1658]  = 255;
  ram[1659]  = 255;
  ram[1660]  = 255;
  ram[1661]  = 255;
  ram[1662]  = 255;
  ram[1663]  = 255;
  ram[1664]  = 255;
  ram[1665]  = 255;
  ram[1666]  = 255;
  ram[1667]  = 255;
  ram[1668]  = 255;
  ram[1669]  = 255;
  ram[1670]  = 255;
  ram[1671]  = 255;
  ram[1672]  = 255;
  ram[1673]  = 255;
  ram[1674]  = 255;
  ram[1675]  = 255;
  ram[1676]  = 255;
  ram[1677]  = 255;
  ram[1678]  = 255;
  ram[1679]  = 255;
  ram[1680]  = 255;
  ram[1681]  = 255;
  ram[1682]  = 255;
  ram[1683]  = 255;
  ram[1684]  = 255;
  ram[1685]  = 255;
  ram[1686]  = 255;
  ram[1687]  = 255;
  ram[1688]  = 255;
  ram[1689]  = 255;
  ram[1690]  = 255;
  ram[1691]  = 255;
  ram[1692]  = 255;
  ram[1693]  = 255;
  ram[1694]  = 255;
  ram[1695]  = 255;
  ram[1696]  = 255;
  ram[1697]  = 255;
  ram[1698]  = 255;
  ram[1699]  = 255;
  ram[1700]  = 255;
  ram[1701]  = 255;
  ram[1702]  = 255;
  ram[1703]  = 255;
  ram[1704]  = 255;
  ram[1705]  = 255;
  ram[1706]  = 255;
  ram[1707]  = 255;
  ram[1708]  = 255;
  ram[1709]  = 255;
  ram[1710]  = 255;
  ram[1711]  = 255;
  ram[1712]  = 255;
  ram[1713]  = 255;
  ram[1714]  = 255;
  ram[1715]  = 255;
  ram[1716]  = 255;
  ram[1717]  = 255;
  ram[1718]  = 255;
  ram[1719]  = 255;
  ram[1720]  = 255;
  ram[1721]  = 255;
  ram[1722]  = 255;
  ram[1723]  = 255;
  ram[1724]  = 255;
  ram[1725]  = 255;
  ram[1726]  = 255;
  ram[1727]  = 255;
  ram[1728]  = 255;
  ram[1729]  = 255;
  ram[1730]  = 255;
  ram[1731]  = 255;
  ram[1732]  = 255;
  ram[1733]  = 255;
  ram[1734]  = 255;
  ram[1735]  = 255;
  ram[1736]  = 255;
  ram[1737]  = 255;
  ram[1738]  = 255;
  ram[1739]  = 255;
  ram[1740]  = 255;
  ram[1741]  = 255;
  ram[1742]  = 255;
  ram[1743]  = 255;
  ram[1744]  = 255;
  ram[1745]  = 255;
  ram[1746]  = 255;
  ram[1747]  = 255;
  ram[1748]  = 255;
  ram[1749]  = 255;
  ram[1750]  = 255;
  ram[1751]  = 255;
  ram[1752]  = 255;
  ram[1753]  = 255;
  ram[1754]  = 255;
  ram[1755]  = 255;
  ram[1756]  = 255;
  ram[1757]  = 255;
  ram[1758]  = 255;
  ram[1759]  = 255;
  ram[1760]  = 255;
  ram[1761]  = 255;
  ram[1762]  = 255;
  ram[1763]  = 255;
  ram[1764]  = 255;
  ram[1765]  = 255;
  ram[1766]  = 255;
  ram[1767]  = 255;
  ram[1768]  = 255;
  ram[1769]  = 255;
  ram[1770]  = 255;
  ram[1771]  = 255;
  ram[1772]  = 255;
  ram[1773]  = 255;
  ram[1774]  = 255;
  ram[1775]  = 255;
  ram[1776]  = 255;
  ram[1777]  = 255;
  ram[1778]  = 255;
  ram[1779]  = 255;
  ram[1780]  = 255;
  ram[1781]  = 255;
  ram[1782]  = 255;
  ram[1783]  = 255;
  ram[1784]  = 255;
  ram[1785]  = 255;
  ram[1786]  = 255;
  ram[1787]  = 255;
  ram[1788]  = 255;
  ram[1789]  = 255;
  ram[1790]  = 255;
  ram[1791]  = 255;
  ram[1792]  = 255;
  ram[1793]  = 255;
  ram[1794]  = 255;
  ram[1795]  = 255;
  ram[1796]  = 236;
  ram[1797]  = 211;
  ram[1798]  = 243;
  ram[1799]  = 255;
  ram[1800]  = 255;
  ram[1801]  = 234;
  ram[1802]  = 206;
  ram[1803]  = 242;
  ram[1804]  = 255;
  ram[1805]  = 254;
  ram[1806]  = 252;
  ram[1807]  = 255;
  ram[1808]  = 255;
  ram[1809]  = 255;
  ram[1810]  = 255;
  ram[1811]  = 255;
  ram[1812]  = 255;
  ram[1813]  = 255;
  ram[1814]  = 255;
  ram[1815]  = 255;
  ram[1816]  = 255;
  ram[1817]  = 255;
  ram[1818]  = 255;
  ram[1819]  = 255;
  ram[1820]  = 255;
  ram[1821]  = 255;
  ram[1822]  = 255;
  ram[1823]  = 255;
  ram[1824]  = 255;
  ram[1825]  = 255;
  ram[1826]  = 255;
  ram[1827]  = 255;
  ram[1828]  = 255;
  ram[1829]  = 255;
  ram[1830]  = 255;
  ram[1831]  = 255;
  ram[1832]  = 255;
  ram[1833]  = 255;
  ram[1834]  = 255;
  ram[1835]  = 255;
  ram[1836]  = 255;
  ram[1837]  = 255;
  ram[1838]  = 255;
  ram[1839]  = 255;
  ram[1840]  = 255;
  ram[1841]  = 255;
  ram[1842]  = 255;
  ram[1843]  = 255;
  ram[1844]  = 255;
  ram[1845]  = 255;
  ram[1846]  = 255;
  ram[1847]  = 255;
  ram[1848]  = 255;
  ram[1849]  = 255;
  ram[1850]  = 255;
  ram[1851]  = 255;
  ram[1852]  = 255;
  ram[1853]  = 255;
  ram[1854]  = 255;
  ram[1855]  = 255;
  ram[1856]  = 255;
  ram[1857]  = 255;
  ram[1858]  = 255;
  ram[1859]  = 255;
  ram[1860]  = 255;
  ram[1861]  = 255;
  ram[1862]  = 255;
  ram[1863]  = 255;
  ram[1864]  = 255;
  ram[1865]  = 255;
  ram[1866]  = 255;
  ram[1867]  = 255;
  ram[1868]  = 255;
  ram[1869]  = 255;
  ram[1870]  = 255;
  ram[1871]  = 255;
  ram[1872]  = 255;
  ram[1873]  = 255;
  ram[1874]  = 255;
  ram[1875]  = 255;
  ram[1876]  = 255;
  ram[1877]  = 255;
  ram[1878]  = 255;
  ram[1879]  = 255;
  ram[1880]  = 255;
  ram[1881]  = 255;
  ram[1882]  = 255;
  ram[1883]  = 255;
  ram[1884]  = 255;
  ram[1885]  = 255;
  ram[1886]  = 255;
  ram[1887]  = 255;
  ram[1888]  = 255;
  ram[1889]  = 255;
  ram[1890]  = 255;
  ram[1891]  = 255;
  ram[1892]  = 255;
  ram[1893]  = 255;
  ram[1894]  = 255;
  ram[1895]  = 255;
  ram[1896]  = 255;
  ram[1897]  = 255;
  ram[1898]  = 255;
  ram[1899]  = 255;
  ram[1900]  = 255;
  ram[1901]  = 255;
  ram[1902]  = 255;
  ram[1903]  = 255;
  ram[1904]  = 255;
  ram[1905]  = 255;
  ram[1906]  = 255;
  ram[1907]  = 255;
  ram[1908]  = 255;
  ram[1909]  = 255;
  ram[1910]  = 255;
  ram[1911]  = 255;
  ram[1912]  = 255;
  ram[1913]  = 255;
  ram[1914]  = 255;
  ram[1915]  = 255;
  ram[1916]  = 255;
  ram[1917]  = 255;
  ram[1918]  = 255;
  ram[1919]  = 255;
  ram[1920]  = 255;
  ram[1921]  = 255;
  ram[1922]  = 255;
  ram[1923]  = 255;
  ram[1924]  = 255;
  ram[1925]  = 255;
  ram[1926]  = 255;
  ram[1927]  = 255;
  ram[1928]  = 255;
  ram[1929]  = 255;
  ram[1930]  = 255;
  ram[1931]  = 255;
  ram[1932]  = 255;
  ram[1933]  = 255;
  ram[1934]  = 255;
  ram[1935]  = 255;
  ram[1936]  = 255;
  ram[1937]  = 255;
  ram[1938]  = 255;
  ram[1939]  = 255;
  ram[1940]  = 255;
  ram[1941]  = 255;
  ram[1942]  = 255;
  ram[1943]  = 255;
  ram[1944]  = 255;
  ram[1945]  = 255;
  ram[1946]  = 255;
  ram[1947]  = 255;
  ram[1948]  = 255;
  ram[1949]  = 255;
  ram[1950]  = 255;
  ram[1951]  = 255;
  ram[1952]  = 255;
  ram[1953]  = 255;
  ram[1954]  = 255;
  ram[1955]  = 255;
  ram[1956]  = 255;
  ram[1957]  = 255;
  ram[1958]  = 255;
  ram[1959]  = 255;
  ram[1960]  = 255;
  ram[1961]  = 255;
  ram[1962]  = 255;
  ram[1963]  = 255;
  ram[1964]  = 255;
  ram[1965]  = 255;
  ram[1966]  = 255;
  ram[1967]  = 255;
  ram[1968]  = 255;
  ram[1969]  = 255;
  ram[1970]  = 255;
  ram[1971]  = 255;
  ram[1972]  = 255;
  ram[1973]  = 255;
  ram[1974]  = 255;
  ram[1975]  = 255;
  ram[1976]  = 255;
  ram[1977]  = 255;
  ram[1978]  = 255;
  ram[1979]  = 255;
  ram[1980]  = 255;
  ram[1981]  = 255;
  ram[1982]  = 255;
  ram[1983]  = 255;
  ram[1984]  = 255;
  ram[1985]  = 255;
  ram[1986]  = 255;
  ram[1987]  = 255;
  ram[1988]  = 255;
  ram[1989]  = 255;
  ram[1990]  = 255;
  ram[1991]  = 255;
  ram[1992]  = 255;
  ram[1993]  = 255;
  ram[1994]  = 255;
  ram[1995]  = 255;
  ram[1996]  = 236;
  ram[1997]  = 211;
  ram[1998]  = 243;
  ram[1999]  = 255;
  ram[2000]  = 255;
  ram[2001]  = 234;
  ram[2002]  = 206;
  ram[2003]  = 242;
  ram[2004]  = 255;
  ram[2005]  = 254;
  ram[2006]  = 252;
  ram[2007]  = 255;
  ram[2008]  = 255;
  ram[2009]  = 255;
  ram[2010]  = 255;
  ram[2011]  = 255;
  ram[2012]  = 255;
  ram[2013]  = 255;
  ram[2014]  = 255;
  ram[2015]  = 255;
  ram[2016]  = 255;
  ram[2017]  = 255;
  ram[2018]  = 255;
  ram[2019]  = 255;
  ram[2020]  = 255;
  ram[2021]  = 255;
  ram[2022]  = 255;
  ram[2023]  = 255;
  ram[2024]  = 255;
  ram[2025]  = 255;
  ram[2026]  = 255;
  ram[2027]  = 255;
  ram[2028]  = 255;
  ram[2029]  = 255;
  ram[2030]  = 255;
  ram[2031]  = 255;
  ram[2032]  = 255;
  ram[2033]  = 255;
  ram[2034]  = 255;
  ram[2035]  = 255;
  ram[2036]  = 255;
  ram[2037]  = 255;
  ram[2038]  = 255;
  ram[2039]  = 255;
  ram[2040]  = 255;
  ram[2041]  = 255;
  ram[2042]  = 255;
  ram[2043]  = 255;
  ram[2044]  = 255;
  ram[2045]  = 255;
  ram[2046]  = 255;
  ram[2047]  = 255;
  ram[2048]  = 255;
  ram[2049]  = 255;
  ram[2050]  = 255;
  ram[2051]  = 255;
  ram[2052]  = 255;
  ram[2053]  = 255;
  ram[2054]  = 255;
  ram[2055]  = 255;
  ram[2056]  = 255;
  ram[2057]  = 255;
  ram[2058]  = 255;
  ram[2059]  = 255;
  ram[2060]  = 255;
  ram[2061]  = 255;
  ram[2062]  = 255;
  ram[2063]  = 255;
  ram[2064]  = 255;
  ram[2065]  = 255;
  ram[2066]  = 255;
  ram[2067]  = 255;
  ram[2068]  = 255;
  ram[2069]  = 255;
  ram[2070]  = 255;
  ram[2071]  = 255;
  ram[2072]  = 255;
  ram[2073]  = 255;
  ram[2074]  = 255;
  ram[2075]  = 255;
  ram[2076]  = 255;
  ram[2077]  = 255;
  ram[2078]  = 255;
  ram[2079]  = 255;
  ram[2080]  = 255;
  ram[2081]  = 255;
  ram[2082]  = 255;
  ram[2083]  = 255;
  ram[2084]  = 255;
  ram[2085]  = 255;
  ram[2086]  = 255;
  ram[2087]  = 255;
  ram[2088]  = 255;
  ram[2089]  = 255;
  ram[2090]  = 255;
  ram[2091]  = 255;
  ram[2092]  = 255;
  ram[2093]  = 255;
  ram[2094]  = 255;
  ram[2095]  = 255;
  ram[2096]  = 255;
  ram[2097]  = 255;
  ram[2098]  = 255;
  ram[2099]  = 255;
  ram[2100]  = 255;
  ram[2101]  = 255;
  ram[2102]  = 255;
  ram[2103]  = 255;
  ram[2104]  = 255;
  ram[2105]  = 255;
  ram[2106]  = 255;
  ram[2107]  = 255;
  ram[2108]  = 255;
  ram[2109]  = 255;
  ram[2110]  = 255;
  ram[2111]  = 255;
  ram[2112]  = 255;
  ram[2113]  = 255;
  ram[2114]  = 255;
  ram[2115]  = 255;
  ram[2116]  = 255;
  ram[2117]  = 255;
  ram[2118]  = 255;
  ram[2119]  = 255;
  ram[2120]  = 255;
  ram[2121]  = 255;
  ram[2122]  = 255;
  ram[2123]  = 255;
  ram[2124]  = 255;
  ram[2125]  = 255;
  ram[2126]  = 255;
  ram[2127]  = 255;
  ram[2128]  = 255;
  ram[2129]  = 255;
  ram[2130]  = 255;
  ram[2131]  = 255;
  ram[2132]  = 255;
  ram[2133]  = 255;
  ram[2134]  = 255;
  ram[2135]  = 255;
  ram[2136]  = 255;
  ram[2137]  = 255;
  ram[2138]  = 255;
  ram[2139]  = 255;
  ram[2140]  = 255;
  ram[2141]  = 255;
  ram[2142]  = 255;
  ram[2143]  = 255;
  ram[2144]  = 255;
  ram[2145]  = 255;
  ram[2146]  = 255;
  ram[2147]  = 255;
  ram[2148]  = 255;
  ram[2149]  = 255;
  ram[2150]  = 255;
  ram[2151]  = 255;
  ram[2152]  = 255;
  ram[2153]  = 255;
  ram[2154]  = 255;
  ram[2155]  = 255;
  ram[2156]  = 255;
  ram[2157]  = 255;
  ram[2158]  = 255;
  ram[2159]  = 255;
  ram[2160]  = 255;
  ram[2161]  = 255;
  ram[2162]  = 255;
  ram[2163]  = 255;
  ram[2164]  = 255;
  ram[2165]  = 255;
  ram[2166]  = 255;
  ram[2167]  = 255;
  ram[2168]  = 255;
  ram[2169]  = 255;
  ram[2170]  = 255;
  ram[2171]  = 255;
  ram[2172]  = 255;
  ram[2173]  = 255;
  ram[2174]  = 255;
  ram[2175]  = 255;
  ram[2176]  = 255;
  ram[2177]  = 255;
  ram[2178]  = 255;
  ram[2179]  = 255;
  ram[2180]  = 255;
  ram[2181]  = 255;
  ram[2182]  = 255;
  ram[2183]  = 255;
  ram[2184]  = 255;
  ram[2185]  = 255;
  ram[2186]  = 255;
  ram[2187]  = 255;
  ram[2188]  = 255;
  ram[2189]  = 255;
  ram[2190]  = 255;
  ram[2191]  = 255;
  ram[2192]  = 255;
  ram[2193]  = 255;
  ram[2194]  = 255;
  ram[2195]  = 255;
  ram[2196]  = 236;
  ram[2197]  = 211;
  ram[2198]  = 243;
  ram[2199]  = 255;
  ram[2200]  = 255;
  ram[2201]  = 234;
  ram[2202]  = 207;
  ram[2203]  = 242;
  ram[2204]  = 255;
  ram[2205]  = 254;
  ram[2206]  = 252;
  ram[2207]  = 255;
  ram[2208]  = 255;
  ram[2209]  = 255;
  ram[2210]  = 255;
  ram[2211]  = 255;
  ram[2212]  = 255;
  ram[2213]  = 255;
  ram[2214]  = 255;
  ram[2215]  = 255;
  ram[2216]  = 255;
  ram[2217]  = 255;
  ram[2218]  = 255;
  ram[2219]  = 255;
  ram[2220]  = 255;
  ram[2221]  = 255;
  ram[2222]  = 255;
  ram[2223]  = 255;
  ram[2224]  = 255;
  ram[2225]  = 255;
  ram[2226]  = 255;
  ram[2227]  = 255;
  ram[2228]  = 255;
  ram[2229]  = 255;
  ram[2230]  = 255;
  ram[2231]  = 255;
  ram[2232]  = 255;
  ram[2233]  = 255;
  ram[2234]  = 255;
  ram[2235]  = 255;
  ram[2236]  = 255;
  ram[2237]  = 255;
  ram[2238]  = 255;
  ram[2239]  = 255;
  ram[2240]  = 255;
  ram[2241]  = 255;
  ram[2242]  = 255;
  ram[2243]  = 255;
  ram[2244]  = 255;
  ram[2245]  = 255;
  ram[2246]  = 255;
  ram[2247]  = 255;
  ram[2248]  = 255;
  ram[2249]  = 255;
  ram[2250]  = 255;
  ram[2251]  = 255;
  ram[2252]  = 255;
  ram[2253]  = 255;
  ram[2254]  = 255;
  ram[2255]  = 255;
  ram[2256]  = 255;
  ram[2257]  = 255;
  ram[2258]  = 255;
  ram[2259]  = 255;
  ram[2260]  = 255;
  ram[2261]  = 255;
  ram[2262]  = 255;
  ram[2263]  = 255;
  ram[2264]  = 255;
  ram[2265]  = 255;
  ram[2266]  = 255;
  ram[2267]  = 255;
  ram[2268]  = 255;
  ram[2269]  = 255;
  ram[2270]  = 255;
  ram[2271]  = 255;
  ram[2272]  = 255;
  ram[2273]  = 255;
  ram[2274]  = 255;
  ram[2275]  = 255;
  ram[2276]  = 255;
  ram[2277]  = 255;
  ram[2278]  = 255;
  ram[2279]  = 255;
  ram[2280]  = 255;
  ram[2281]  = 255;
  ram[2282]  = 255;
  ram[2283]  = 255;
  ram[2284]  = 255;
  ram[2285]  = 255;
  ram[2286]  = 255;
  ram[2287]  = 255;
  ram[2288]  = 255;
  ram[2289]  = 255;
  ram[2290]  = 255;
  ram[2291]  = 255;
  ram[2292]  = 255;
  ram[2293]  = 255;
  ram[2294]  = 255;
  ram[2295]  = 255;
  ram[2296]  = 255;
  ram[2297]  = 255;
  ram[2298]  = 255;
  ram[2299]  = 255;
  ram[2300]  = 255;
  ram[2301]  = 255;
  ram[2302]  = 255;
  ram[2303]  = 255;
  ram[2304]  = 255;
  ram[2305]  = 255;
  ram[2306]  = 255;
  ram[2307]  = 255;
  ram[2308]  = 255;
  ram[2309]  = 255;
  ram[2310]  = 255;
  ram[2311]  = 255;
  ram[2312]  = 255;
  ram[2313]  = 255;
  ram[2314]  = 255;
  ram[2315]  = 255;
  ram[2316]  = 255;
  ram[2317]  = 255;
  ram[2318]  = 255;
  ram[2319]  = 255;
  ram[2320]  = 255;
  ram[2321]  = 255;
  ram[2322]  = 255;
  ram[2323]  = 255;
  ram[2324]  = 255;
  ram[2325]  = 255;
  ram[2326]  = 255;
  ram[2327]  = 255;
  ram[2328]  = 255;
  ram[2329]  = 255;
  ram[2330]  = 255;
  ram[2331]  = 255;
  ram[2332]  = 255;
  ram[2333]  = 255;
  ram[2334]  = 255;
  ram[2335]  = 255;
  ram[2336]  = 255;
  ram[2337]  = 255;
  ram[2338]  = 255;
  ram[2339]  = 255;
  ram[2340]  = 255;
  ram[2341]  = 255;
  ram[2342]  = 255;
  ram[2343]  = 255;
  ram[2344]  = 255;
  ram[2345]  = 255;
  ram[2346]  = 255;
  ram[2347]  = 255;
  ram[2348]  = 255;
  ram[2349]  = 255;
  ram[2350]  = 255;
  ram[2351]  = 255;
  ram[2352]  = 255;
  ram[2353]  = 255;
  ram[2354]  = 255;
  ram[2355]  = 255;
  ram[2356]  = 255;
  ram[2357]  = 255;
  ram[2358]  = 255;
  ram[2359]  = 255;
  ram[2360]  = 255;
  ram[2361]  = 255;
  ram[2362]  = 255;
  ram[2363]  = 255;
  ram[2364]  = 255;
  ram[2365]  = 255;
  ram[2366]  = 255;
  ram[2367]  = 255;
  ram[2368]  = 255;
  ram[2369]  = 255;
  ram[2370]  = 255;
  ram[2371]  = 255;
  ram[2372]  = 255;
  ram[2373]  = 255;
  ram[2374]  = 255;
  ram[2375]  = 255;
  ram[2376]  = 255;
  ram[2377]  = 255;
  ram[2378]  = 255;
  ram[2379]  = 255;
  ram[2380]  = 255;
  ram[2381]  = 255;
  ram[2382]  = 255;
  ram[2383]  = 255;
  ram[2384]  = 255;
  ram[2385]  = 255;
  ram[2386]  = 255;
  ram[2387]  = 255;
  ram[2388]  = 255;
  ram[2389]  = 255;
  ram[2390]  = 255;
  ram[2391]  = 255;
  ram[2392]  = 255;
  ram[2393]  = 255;
  ram[2394]  = 255;
  ram[2395]  = 255;
  ram[2396]  = 235;
  ram[2397]  = 211;
  ram[2398]  = 243;
  ram[2399]  = 255;
  ram[2400]  = 253;
  ram[2401]  = 235;
  ram[2402]  = 208;
  ram[2403]  = 242;
  ram[2404]  = 255;
  ram[2405]  = 254;
  ram[2406]  = 252;
  ram[2407]  = 255;
  ram[2408]  = 255;
  ram[2409]  = 255;
  ram[2410]  = 255;
  ram[2411]  = 255;
  ram[2412]  = 255;
  ram[2413]  = 255;
  ram[2414]  = 255;
  ram[2415]  = 255;
  ram[2416]  = 255;
  ram[2417]  = 255;
  ram[2418]  = 255;
  ram[2419]  = 255;
  ram[2420]  = 255;
  ram[2421]  = 255;
  ram[2422]  = 255;
  ram[2423]  = 255;
  ram[2424]  = 255;
  ram[2425]  = 255;
  ram[2426]  = 255;
  ram[2427]  = 255;
  ram[2428]  = 255;
  ram[2429]  = 255;
  ram[2430]  = 255;
  ram[2431]  = 255;
  ram[2432]  = 255;
  ram[2433]  = 255;
  ram[2434]  = 255;
  ram[2435]  = 255;
  ram[2436]  = 255;
  ram[2437]  = 255;
  ram[2438]  = 255;
  ram[2439]  = 255;
  ram[2440]  = 255;
  ram[2441]  = 255;
  ram[2442]  = 255;
  ram[2443]  = 255;
  ram[2444]  = 255;
  ram[2445]  = 255;
  ram[2446]  = 255;
  ram[2447]  = 255;
  ram[2448]  = 255;
  ram[2449]  = 255;
  ram[2450]  = 255;
  ram[2451]  = 255;
  ram[2452]  = 255;
  ram[2453]  = 255;
  ram[2454]  = 255;
  ram[2455]  = 255;
  ram[2456]  = 255;
  ram[2457]  = 255;
  ram[2458]  = 255;
  ram[2459]  = 255;
  ram[2460]  = 255;
  ram[2461]  = 255;
  ram[2462]  = 255;
  ram[2463]  = 255;
  ram[2464]  = 255;
  ram[2465]  = 255;
  ram[2466]  = 255;
  ram[2467]  = 255;
  ram[2468]  = 255;
  ram[2469]  = 255;
  ram[2470]  = 255;
  ram[2471]  = 255;
  ram[2472]  = 255;
  ram[2473]  = 255;
  ram[2474]  = 255;
  ram[2475]  = 255;
  ram[2476]  = 255;
  ram[2477]  = 255;
  ram[2478]  = 255;
  ram[2479]  = 255;
  ram[2480]  = 255;
  ram[2481]  = 255;
  ram[2482]  = 255;
  ram[2483]  = 255;
  ram[2484]  = 255;
  ram[2485]  = 255;
  ram[2486]  = 255;
  ram[2487]  = 255;
  ram[2488]  = 255;
  ram[2489]  = 255;
  ram[2490]  = 255;
  ram[2491]  = 255;
  ram[2492]  = 255;
  ram[2493]  = 255;
  ram[2494]  = 255;
  ram[2495]  = 255;
  ram[2496]  = 255;
  ram[2497]  = 255;
  ram[2498]  = 255;
  ram[2499]  = 255;
  ram[2500]  = 255;
  ram[2501]  = 255;
  ram[2502]  = 255;
  ram[2503]  = 255;
  ram[2504]  = 255;
  ram[2505]  = 255;
  ram[2506]  = 255;
  ram[2507]  = 255;
  ram[2508]  = 255;
  ram[2509]  = 255;
  ram[2510]  = 255;
  ram[2511]  = 255;
  ram[2512]  = 255;
  ram[2513]  = 255;
  ram[2514]  = 255;
  ram[2515]  = 255;
  ram[2516]  = 255;
  ram[2517]  = 255;
  ram[2518]  = 255;
  ram[2519]  = 255;
  ram[2520]  = 255;
  ram[2521]  = 255;
  ram[2522]  = 255;
  ram[2523]  = 255;
  ram[2524]  = 255;
  ram[2525]  = 255;
  ram[2526]  = 255;
  ram[2527]  = 255;
  ram[2528]  = 255;
  ram[2529]  = 255;
  ram[2530]  = 255;
  ram[2531]  = 255;
  ram[2532]  = 255;
  ram[2533]  = 255;
  ram[2534]  = 255;
  ram[2535]  = 255;
  ram[2536]  = 255;
  ram[2537]  = 255;
  ram[2538]  = 255;
  ram[2539]  = 255;
  ram[2540]  = 255;
  ram[2541]  = 255;
  ram[2542]  = 255;
  ram[2543]  = 255;
  ram[2544]  = 255;
  ram[2545]  = 255;
  ram[2546]  = 255;
  ram[2547]  = 255;
  ram[2548]  = 255;
  ram[2549]  = 255;
  ram[2550]  = 255;
  ram[2551]  = 255;
  ram[2552]  = 255;
  ram[2553]  = 255;
  ram[2554]  = 255;
  ram[2555]  = 255;
  ram[2556]  = 255;
  ram[2557]  = 255;
  ram[2558]  = 255;
  ram[2559]  = 255;
  ram[2560]  = 255;
  ram[2561]  = 255;
  ram[2562]  = 255;
  ram[2563]  = 255;
  ram[2564]  = 255;
  ram[2565]  = 255;
  ram[2566]  = 255;
  ram[2567]  = 255;
  ram[2568]  = 255;
  ram[2569]  = 255;
  ram[2570]  = 255;
  ram[2571]  = 255;
  ram[2572]  = 255;
  ram[2573]  = 255;
  ram[2574]  = 255;
  ram[2575]  = 255;
  ram[2576]  = 255;
  ram[2577]  = 255;
  ram[2578]  = 255;
  ram[2579]  = 255;
  ram[2580]  = 255;
  ram[2581]  = 255;
  ram[2582]  = 255;
  ram[2583]  = 255;
  ram[2584]  = 255;
  ram[2585]  = 255;
  ram[2586]  = 255;
  ram[2587]  = 255;
  ram[2588]  = 255;
  ram[2589]  = 255;
  ram[2590]  = 255;
  ram[2591]  = 255;
  ram[2592]  = 255;
  ram[2593]  = 255;
  ram[2594]  = 255;
  ram[2595]  = 255;
  ram[2596]  = 235;
  ram[2597]  = 212;
  ram[2598]  = 243;
  ram[2599]  = 255;
  ram[2600]  = 252;
  ram[2601]  = 235;
  ram[2602]  = 209;
  ram[2603]  = 242;
  ram[2604]  = 255;
  ram[2605]  = 254;
  ram[2606]  = 252;
  ram[2607]  = 255;
  ram[2608]  = 255;
  ram[2609]  = 255;
  ram[2610]  = 255;
  ram[2611]  = 255;
  ram[2612]  = 255;
  ram[2613]  = 255;
  ram[2614]  = 255;
  ram[2615]  = 255;
  ram[2616]  = 255;
  ram[2617]  = 255;
  ram[2618]  = 255;
  ram[2619]  = 255;
  ram[2620]  = 255;
  ram[2621]  = 255;
  ram[2622]  = 255;
  ram[2623]  = 255;
  ram[2624]  = 255;
  ram[2625]  = 255;
  ram[2626]  = 255;
  ram[2627]  = 255;
  ram[2628]  = 255;
  ram[2629]  = 255;
  ram[2630]  = 255;
  ram[2631]  = 255;
  ram[2632]  = 255;
  ram[2633]  = 255;
  ram[2634]  = 255;
  ram[2635]  = 255;
  ram[2636]  = 255;
  ram[2637]  = 255;
  ram[2638]  = 255;
  ram[2639]  = 255;
  ram[2640]  = 255;
  ram[2641]  = 255;
  ram[2642]  = 255;
  ram[2643]  = 255;
  ram[2644]  = 255;
  ram[2645]  = 255;
  ram[2646]  = 255;
  ram[2647]  = 255;
  ram[2648]  = 255;
  ram[2649]  = 255;
  ram[2650]  = 255;
  ram[2651]  = 255;
  ram[2652]  = 255;
  ram[2653]  = 255;
  ram[2654]  = 255;
  ram[2655]  = 255;
  ram[2656]  = 255;
  ram[2657]  = 255;
  ram[2658]  = 255;
  ram[2659]  = 255;
  ram[2660]  = 255;
  ram[2661]  = 255;
  ram[2662]  = 255;
  ram[2663]  = 255;
  ram[2664]  = 255;
  ram[2665]  = 255;
  ram[2666]  = 255;
  ram[2667]  = 255;
  ram[2668]  = 255;
  ram[2669]  = 255;
  ram[2670]  = 255;
  ram[2671]  = 255;
  ram[2672]  = 255;
  ram[2673]  = 255;
  ram[2674]  = 255;
  ram[2675]  = 255;
  ram[2676]  = 255;
  ram[2677]  = 255;
  ram[2678]  = 255;
  ram[2679]  = 255;
  ram[2680]  = 255;
  ram[2681]  = 255;
  ram[2682]  = 255;
  ram[2683]  = 255;
  ram[2684]  = 255;
  ram[2685]  = 255;
  ram[2686]  = 255;
  ram[2687]  = 255;
  ram[2688]  = 255;
  ram[2689]  = 255;
  ram[2690]  = 255;
  ram[2691]  = 255;
  ram[2692]  = 255;
  ram[2693]  = 255;
  ram[2694]  = 255;
  ram[2695]  = 255;
  ram[2696]  = 255;
  ram[2697]  = 255;
  ram[2698]  = 255;
  ram[2699]  = 255;
  ram[2700]  = 255;
  ram[2701]  = 255;
  ram[2702]  = 255;
  ram[2703]  = 255;
  ram[2704]  = 255;
  ram[2705]  = 255;
  ram[2706]  = 255;
  ram[2707]  = 255;
  ram[2708]  = 255;
  ram[2709]  = 255;
  ram[2710]  = 255;
  ram[2711]  = 255;
  ram[2712]  = 255;
  ram[2713]  = 255;
  ram[2714]  = 255;
  ram[2715]  = 255;
  ram[2716]  = 255;
  ram[2717]  = 255;
  ram[2718]  = 255;
  ram[2719]  = 255;
  ram[2720]  = 255;
  ram[2721]  = 255;
  ram[2722]  = 255;
  ram[2723]  = 255;
  ram[2724]  = 255;
  ram[2725]  = 255;
  ram[2726]  = 255;
  ram[2727]  = 255;
  ram[2728]  = 255;
  ram[2729]  = 255;
  ram[2730]  = 255;
  ram[2731]  = 255;
  ram[2732]  = 255;
  ram[2733]  = 255;
  ram[2734]  = 255;
  ram[2735]  = 255;
  ram[2736]  = 255;
  ram[2737]  = 255;
  ram[2738]  = 255;
  ram[2739]  = 255;
  ram[2740]  = 255;
  ram[2741]  = 255;
  ram[2742]  = 255;
  ram[2743]  = 255;
  ram[2744]  = 255;
  ram[2745]  = 255;
  ram[2746]  = 255;
  ram[2747]  = 255;
  ram[2748]  = 255;
  ram[2749]  = 255;
  ram[2750]  = 255;
  ram[2751]  = 255;
  ram[2752]  = 255;
  ram[2753]  = 255;
  ram[2754]  = 255;
  ram[2755]  = 255;
  ram[2756]  = 255;
  ram[2757]  = 255;
  ram[2758]  = 255;
  ram[2759]  = 255;
  ram[2760]  = 255;
  ram[2761]  = 255;
  ram[2762]  = 255;
  ram[2763]  = 255;
  ram[2764]  = 255;
  ram[2765]  = 255;
  ram[2766]  = 255;
  ram[2767]  = 255;
  ram[2768]  = 255;
  ram[2769]  = 255;
  ram[2770]  = 255;
  ram[2771]  = 255;
  ram[2772]  = 255;
  ram[2773]  = 255;
  ram[2774]  = 255;
  ram[2775]  = 255;
  ram[2776]  = 255;
  ram[2777]  = 255;
  ram[2778]  = 255;
  ram[2779]  = 255;
  ram[2780]  = 255;
  ram[2781]  = 255;
  ram[2782]  = 255;
  ram[2783]  = 255;
  ram[2784]  = 255;
  ram[2785]  = 255;
  ram[2786]  = 255;
  ram[2787]  = 255;
  ram[2788]  = 255;
  ram[2789]  = 255;
  ram[2790]  = 255;
  ram[2791]  = 255;
  ram[2792]  = 255;
  ram[2793]  = 255;
  ram[2794]  = 255;
  ram[2795]  = 255;
  ram[2796]  = 236;
  ram[2797]  = 211;
  ram[2798]  = 243;
  ram[2799]  = 255;
  ram[2800]  = 253;
  ram[2801]  = 235;
  ram[2802]  = 209;
  ram[2803]  = 242;
  ram[2804]  = 255;
  ram[2805]  = 254;
  ram[2806]  = 252;
  ram[2807]  = 255;
  ram[2808]  = 255;
  ram[2809]  = 255;
  ram[2810]  = 255;
  ram[2811]  = 255;
  ram[2812]  = 255;
  ram[2813]  = 255;
  ram[2814]  = 255;
  ram[2815]  = 255;
  ram[2816]  = 255;
  ram[2817]  = 255;
  ram[2818]  = 255;
  ram[2819]  = 255;
  ram[2820]  = 255;
  ram[2821]  = 255;
  ram[2822]  = 255;
  ram[2823]  = 255;
  ram[2824]  = 255;
  ram[2825]  = 255;
  ram[2826]  = 255;
  ram[2827]  = 255;
  ram[2828]  = 255;
  ram[2829]  = 255;
  ram[2830]  = 255;
  ram[2831]  = 255;
  ram[2832]  = 255;
  ram[2833]  = 255;
  ram[2834]  = 255;
  ram[2835]  = 255;
  ram[2836]  = 255;
  ram[2837]  = 255;
  ram[2838]  = 255;
  ram[2839]  = 255;
  ram[2840]  = 255;
  ram[2841]  = 255;
  ram[2842]  = 255;
  ram[2843]  = 255;
  ram[2844]  = 255;
  ram[2845]  = 255;
  ram[2846]  = 255;
  ram[2847]  = 255;
  ram[2848]  = 255;
  ram[2849]  = 255;
  ram[2850]  = 255;
  ram[2851]  = 255;
  ram[2852]  = 255;
  ram[2853]  = 255;
  ram[2854]  = 255;
  ram[2855]  = 255;
  ram[2856]  = 255;
  ram[2857]  = 255;
  ram[2858]  = 255;
  ram[2859]  = 255;
  ram[2860]  = 255;
  ram[2861]  = 255;
  ram[2862]  = 255;
  ram[2863]  = 255;
  ram[2864]  = 255;
  ram[2865]  = 255;
  ram[2866]  = 255;
  ram[2867]  = 255;
  ram[2868]  = 255;
  ram[2869]  = 255;
  ram[2870]  = 255;
  ram[2871]  = 255;
  ram[2872]  = 255;
  ram[2873]  = 255;
  ram[2874]  = 255;
  ram[2875]  = 255;
  ram[2876]  = 255;
  ram[2877]  = 255;
  ram[2878]  = 255;
  ram[2879]  = 255;
  ram[2880]  = 255;
  ram[2881]  = 255;
  ram[2882]  = 255;
  ram[2883]  = 255;
  ram[2884]  = 255;
  ram[2885]  = 255;
  ram[2886]  = 255;
  ram[2887]  = 255;
  ram[2888]  = 255;
  ram[2889]  = 255;
  ram[2890]  = 255;
  ram[2891]  = 255;
  ram[2892]  = 255;
  ram[2893]  = 255;
  ram[2894]  = 255;
  ram[2895]  = 255;
  ram[2896]  = 255;
  ram[2897]  = 255;
  ram[2898]  = 255;
  ram[2899]  = 255;
  ram[2900]  = 255;
  ram[2901]  = 255;
  ram[2902]  = 255;
  ram[2903]  = 255;
  ram[2904]  = 255;
  ram[2905]  = 255;
  ram[2906]  = 255;
  ram[2907]  = 255;
  ram[2908]  = 255;
  ram[2909]  = 255;
  ram[2910]  = 255;
  ram[2911]  = 255;
  ram[2912]  = 255;
  ram[2913]  = 255;
  ram[2914]  = 255;
  ram[2915]  = 255;
  ram[2916]  = 255;
  ram[2917]  = 255;
  ram[2918]  = 255;
  ram[2919]  = 255;
  ram[2920]  = 255;
  ram[2921]  = 255;
  ram[2922]  = 255;
  ram[2923]  = 255;
  ram[2924]  = 255;
  ram[2925]  = 255;
  ram[2926]  = 255;
  ram[2927]  = 255;
  ram[2928]  = 255;
  ram[2929]  = 255;
  ram[2930]  = 255;
  ram[2931]  = 255;
  ram[2932]  = 255;
  ram[2933]  = 255;
  ram[2934]  = 255;
  ram[2935]  = 255;
  ram[2936]  = 255;
  ram[2937]  = 255;
  ram[2938]  = 255;
  ram[2939]  = 255;
  ram[2940]  = 255;
  ram[2941]  = 255;
  ram[2942]  = 255;
  ram[2943]  = 255;
  ram[2944]  = 255;
  ram[2945]  = 255;
  ram[2946]  = 255;
  ram[2947]  = 255;
  ram[2948]  = 255;
  ram[2949]  = 255;
  ram[2950]  = 255;
  ram[2951]  = 255;
  ram[2952]  = 255;
  ram[2953]  = 255;
  ram[2954]  = 255;
  ram[2955]  = 255;
  ram[2956]  = 255;
  ram[2957]  = 255;
  ram[2958]  = 255;
  ram[2959]  = 255;
  ram[2960]  = 255;
  ram[2961]  = 255;
  ram[2962]  = 255;
  ram[2963]  = 255;
  ram[2964]  = 255;
  ram[2965]  = 255;
  ram[2966]  = 255;
  ram[2967]  = 255;
  ram[2968]  = 255;
  ram[2969]  = 255;
  ram[2970]  = 255;
  ram[2971]  = 255;
  ram[2972]  = 255;
  ram[2973]  = 255;
  ram[2974]  = 255;
  ram[2975]  = 255;
  ram[2976]  = 255;
  ram[2977]  = 255;
  ram[2978]  = 255;
  ram[2979]  = 255;
  ram[2980]  = 255;
  ram[2981]  = 255;
  ram[2982]  = 255;
  ram[2983]  = 255;
  ram[2984]  = 255;
  ram[2985]  = 255;
  ram[2986]  = 255;
  ram[2987]  = 255;
  ram[2988]  = 255;
  ram[2989]  = 255;
  ram[2990]  = 255;
  ram[2991]  = 255;
  ram[2992]  = 255;
  ram[2993]  = 255;
  ram[2994]  = 255;
  ram[2995]  = 255;
  ram[2996]  = 236;
  ram[2997]  = 211;
  ram[2998]  = 243;
  ram[2999]  = 255;
  ram[3000]  = 253;
  ram[3001]  = 235;
  ram[3002]  = 209;
  ram[3003]  = 242;
  ram[3004]  = 255;
  ram[3005]  = 254;
  ram[3006]  = 252;
  ram[3007]  = 255;
  ram[3008]  = 255;
  ram[3009]  = 255;
  ram[3010]  = 255;
  ram[3011]  = 255;
  ram[3012]  = 255;
  ram[3013]  = 255;
  ram[3014]  = 254;
  ram[3015]  = 253;
  ram[3016]  = 252;
  ram[3017]  = 255;
  ram[3018]  = 255;
  ram[3019]  = 254;
  ram[3020]  = 254;
  ram[3021]  = 253;
  ram[3022]  = 254;
  ram[3023]  = 252;
  ram[3024]  = 253;
  ram[3025]  = 255;
  ram[3026]  = 255;
  ram[3027]  = 255;
  ram[3028]  = 255;
  ram[3029]  = 255;
  ram[3030]  = 255;
  ram[3031]  = 255;
  ram[3032]  = 255;
  ram[3033]  = 255;
  ram[3034]  = 255;
  ram[3035]  = 255;
  ram[3036]  = 255;
  ram[3037]  = 255;
  ram[3038]  = 255;
  ram[3039]  = 255;
  ram[3040]  = 255;
  ram[3041]  = 255;
  ram[3042]  = 255;
  ram[3043]  = 255;
  ram[3044]  = 255;
  ram[3045]  = 255;
  ram[3046]  = 255;
  ram[3047]  = 255;
  ram[3048]  = 255;
  ram[3049]  = 255;
  ram[3050]  = 255;
  ram[3051]  = 255;
  ram[3052]  = 255;
  ram[3053]  = 255;
  ram[3054]  = 255;
  ram[3055]  = 255;
  ram[3056]  = 255;
  ram[3057]  = 255;
  ram[3058]  = 255;
  ram[3059]  = 255;
  ram[3060]  = 255;
  ram[3061]  = 254;
  ram[3062]  = 253;
  ram[3063]  = 255;
  ram[3064]  = 255;
  ram[3065]  = 254;
  ram[3066]  = 255;
  ram[3067]  = 255;
  ram[3068]  = 255;
  ram[3069]  = 255;
  ram[3070]  = 255;
  ram[3071]  = 255;
  ram[3072]  = 255;
  ram[3073]  = 255;
  ram[3074]  = 255;
  ram[3075]  = 255;
  ram[3076]  = 255;
  ram[3077]  = 255;
  ram[3078]  = 255;
  ram[3079]  = 255;
  ram[3080]  = 255;
  ram[3081]  = 255;
  ram[3082]  = 255;
  ram[3083]  = 255;
  ram[3084]  = 254;
  ram[3085]  = 255;
  ram[3086]  = 255;
  ram[3087]  = 255;
  ram[3088]  = 255;
  ram[3089]  = 255;
  ram[3090]  = 255;
  ram[3091]  = 255;
  ram[3092]  = 255;
  ram[3093]  = 255;
  ram[3094]  = 255;
  ram[3095]  = 255;
  ram[3096]  = 255;
  ram[3097]  = 255;
  ram[3098]  = 255;
  ram[3099]  = 255;
  ram[3100]  = 255;
  ram[3101]  = 255;
  ram[3102]  = 255;
  ram[3103]  = 255;
  ram[3104]  = 255;
  ram[3105]  = 255;
  ram[3106]  = 255;
  ram[3107]  = 255;
  ram[3108]  = 255;
  ram[3109]  = 255;
  ram[3110]  = 255;
  ram[3111]  = 255;
  ram[3112]  = 255;
  ram[3113]  = 255;
  ram[3114]  = 255;
  ram[3115]  = 255;
  ram[3116]  = 255;
  ram[3117]  = 255;
  ram[3118]  = 255;
  ram[3119]  = 255;
  ram[3120]  = 255;
  ram[3121]  = 255;
  ram[3122]  = 255;
  ram[3123]  = 255;
  ram[3124]  = 255;
  ram[3125]  = 255;
  ram[3126]  = 255;
  ram[3127]  = 255;
  ram[3128]  = 255;
  ram[3129]  = 255;
  ram[3130]  = 255;
  ram[3131]  = 255;
  ram[3132]  = 255;
  ram[3133]  = 255;
  ram[3134]  = 255;
  ram[3135]  = 255;
  ram[3136]  = 255;
  ram[3137]  = 255;
  ram[3138]  = 255;
  ram[3139]  = 255;
  ram[3140]  = 255;
  ram[3141]  = 255;
  ram[3142]  = 255;
  ram[3143]  = 255;
  ram[3144]  = 255;
  ram[3145]  = 255;
  ram[3146]  = 255;
  ram[3147]  = 255;
  ram[3148]  = 255;
  ram[3149]  = 255;
  ram[3150]  = 255;
  ram[3151]  = 255;
  ram[3152]  = 255;
  ram[3153]  = 255;
  ram[3154]  = 255;
  ram[3155]  = 255;
  ram[3156]  = 255;
  ram[3157]  = 255;
  ram[3158]  = 255;
  ram[3159]  = 255;
  ram[3160]  = 255;
  ram[3161]  = 255;
  ram[3162]  = 255;
  ram[3163]  = 255;
  ram[3164]  = 255;
  ram[3165]  = 255;
  ram[3166]  = 255;
  ram[3167]  = 255;
  ram[3168]  = 255;
  ram[3169]  = 255;
  ram[3170]  = 255;
  ram[3171]  = 255;
  ram[3172]  = 255;
  ram[3173]  = 255;
  ram[3174]  = 255;
  ram[3175]  = 255;
  ram[3176]  = 255;
  ram[3177]  = 255;
  ram[3178]  = 255;
  ram[3179]  = 255;
  ram[3180]  = 255;
  ram[3181]  = 255;
  ram[3182]  = 255;
  ram[3183]  = 255;
  ram[3184]  = 255;
  ram[3185]  = 255;
  ram[3186]  = 255;
  ram[3187]  = 255;
  ram[3188]  = 255;
  ram[3189]  = 255;
  ram[3190]  = 255;
  ram[3191]  = 255;
  ram[3192]  = 255;
  ram[3193]  = 255;
  ram[3194]  = 255;
  ram[3195]  = 255;
  ram[3196]  = 236;
  ram[3197]  = 211;
  ram[3198]  = 243;
  ram[3199]  = 255;
  ram[3200]  = 253;
  ram[3201]  = 235;
  ram[3202]  = 209;
  ram[3203]  = 242;
  ram[3204]  = 255;
  ram[3205]  = 254;
  ram[3206]  = 252;
  ram[3207]  = 255;
  ram[3208]  = 255;
  ram[3209]  = 255;
  ram[3210]  = 255;
  ram[3211]  = 255;
  ram[3212]  = 255;
  ram[3213]  = 255;
  ram[3214]  = 254;
  ram[3215]  = 251;
  ram[3216]  = 253;
  ram[3217]  = 255;
  ram[3218]  = 255;
  ram[3219]  = 255;
  ram[3220]  = 255;
  ram[3221]  = 255;
  ram[3222]  = 251;
  ram[3223]  = 253;
  ram[3224]  = 254;
  ram[3225]  = 255;
  ram[3226]  = 255;
  ram[3227]  = 255;
  ram[3228]  = 255;
  ram[3229]  = 255;
  ram[3230]  = 255;
  ram[3231]  = 255;
  ram[3232]  = 255;
  ram[3233]  = 255;
  ram[3234]  = 255;
  ram[3235]  = 255;
  ram[3236]  = 255;
  ram[3237]  = 255;
  ram[3238]  = 255;
  ram[3239]  = 255;
  ram[3240]  = 255;
  ram[3241]  = 255;
  ram[3242]  = 255;
  ram[3243]  = 255;
  ram[3244]  = 255;
  ram[3245]  = 255;
  ram[3246]  = 255;
  ram[3247]  = 255;
  ram[3248]  = 255;
  ram[3249]  = 255;
  ram[3250]  = 255;
  ram[3251]  = 255;
  ram[3252]  = 255;
  ram[3253]  = 255;
  ram[3254]  = 255;
  ram[3255]  = 255;
  ram[3256]  = 255;
  ram[3257]  = 255;
  ram[3258]  = 255;
  ram[3259]  = 255;
  ram[3260]  = 255;
  ram[3261]  = 253;
  ram[3262]  = 255;
  ram[3263]  = 229;
  ram[3264]  = 200;
  ram[3265]  = 255;
  ram[3266]  = 254;
  ram[3267]  = 255;
  ram[3268]  = 255;
  ram[3269]  = 255;
  ram[3270]  = 255;
  ram[3271]  = 255;
  ram[3272]  = 255;
  ram[3273]  = 255;
  ram[3274]  = 255;
  ram[3275]  = 255;
  ram[3276]  = 255;
  ram[3277]  = 255;
  ram[3278]  = 255;
  ram[3279]  = 255;
  ram[3280]  = 255;
  ram[3281]  = 255;
  ram[3282]  = 255;
  ram[3283]  = 255;
  ram[3284]  = 255;
  ram[3285]  = 235;
  ram[3286]  = 200;
  ram[3287]  = 254;
  ram[3288]  = 253;
  ram[3289]  = 255;
  ram[3290]  = 255;
  ram[3291]  = 255;
  ram[3292]  = 255;
  ram[3293]  = 255;
  ram[3294]  = 255;
  ram[3295]  = 255;
  ram[3296]  = 255;
  ram[3297]  = 255;
  ram[3298]  = 255;
  ram[3299]  = 255;
  ram[3300]  = 255;
  ram[3301]  = 255;
  ram[3302]  = 255;
  ram[3303]  = 255;
  ram[3304]  = 255;
  ram[3305]  = 255;
  ram[3306]  = 255;
  ram[3307]  = 255;
  ram[3308]  = 255;
  ram[3309]  = 255;
  ram[3310]  = 255;
  ram[3311]  = 255;
  ram[3312]  = 255;
  ram[3313]  = 255;
  ram[3314]  = 255;
  ram[3315]  = 255;
  ram[3316]  = 255;
  ram[3317]  = 255;
  ram[3318]  = 255;
  ram[3319]  = 255;
  ram[3320]  = 255;
  ram[3321]  = 255;
  ram[3322]  = 255;
  ram[3323]  = 255;
  ram[3324]  = 255;
  ram[3325]  = 255;
  ram[3326]  = 255;
  ram[3327]  = 255;
  ram[3328]  = 255;
  ram[3329]  = 255;
  ram[3330]  = 255;
  ram[3331]  = 255;
  ram[3332]  = 255;
  ram[3333]  = 255;
  ram[3334]  = 255;
  ram[3335]  = 255;
  ram[3336]  = 255;
  ram[3337]  = 255;
  ram[3338]  = 255;
  ram[3339]  = 255;
  ram[3340]  = 255;
  ram[3341]  = 255;
  ram[3342]  = 255;
  ram[3343]  = 255;
  ram[3344]  = 255;
  ram[3345]  = 255;
  ram[3346]  = 255;
  ram[3347]  = 255;
  ram[3348]  = 255;
  ram[3349]  = 255;
  ram[3350]  = 255;
  ram[3351]  = 255;
  ram[3352]  = 255;
  ram[3353]  = 255;
  ram[3354]  = 255;
  ram[3355]  = 255;
  ram[3356]  = 255;
  ram[3357]  = 255;
  ram[3358]  = 255;
  ram[3359]  = 255;
  ram[3360]  = 255;
  ram[3361]  = 255;
  ram[3362]  = 255;
  ram[3363]  = 255;
  ram[3364]  = 255;
  ram[3365]  = 255;
  ram[3366]  = 255;
  ram[3367]  = 255;
  ram[3368]  = 255;
  ram[3369]  = 255;
  ram[3370]  = 255;
  ram[3371]  = 255;
  ram[3372]  = 255;
  ram[3373]  = 255;
  ram[3374]  = 255;
  ram[3375]  = 255;
  ram[3376]  = 255;
  ram[3377]  = 255;
  ram[3378]  = 255;
  ram[3379]  = 255;
  ram[3380]  = 255;
  ram[3381]  = 255;
  ram[3382]  = 255;
  ram[3383]  = 255;
  ram[3384]  = 255;
  ram[3385]  = 255;
  ram[3386]  = 255;
  ram[3387]  = 255;
  ram[3388]  = 255;
  ram[3389]  = 255;
  ram[3390]  = 255;
  ram[3391]  = 255;
  ram[3392]  = 255;
  ram[3393]  = 255;
  ram[3394]  = 255;
  ram[3395]  = 255;
  ram[3396]  = 236;
  ram[3397]  = 211;
  ram[3398]  = 243;
  ram[3399]  = 255;
  ram[3400]  = 253;
  ram[3401]  = 235;
  ram[3402]  = 209;
  ram[3403]  = 242;
  ram[3404]  = 255;
  ram[3405]  = 254;
  ram[3406]  = 252;
  ram[3407]  = 255;
  ram[3408]  = 255;
  ram[3409]  = 255;
  ram[3410]  = 255;
  ram[3411]  = 255;
  ram[3412]  = 255;
  ram[3413]  = 255;
  ram[3414]  = 254;
  ram[3415]  = 255;
  ram[3416]  = 225;
  ram[3417]  = 158;
  ram[3418]  = 166;
  ram[3419]  = 166;
  ram[3420]  = 170;
  ram[3421]  = 225;
  ram[3422]  = 255;
  ram[3423]  = 253;
  ram[3424]  = 254;
  ram[3425]  = 255;
  ram[3426]  = 255;
  ram[3427]  = 255;
  ram[3428]  = 255;
  ram[3429]  = 255;
  ram[3430]  = 255;
  ram[3431]  = 255;
  ram[3432]  = 255;
  ram[3433]  = 255;
  ram[3434]  = 255;
  ram[3435]  = 255;
  ram[3436]  = 255;
  ram[3437]  = 255;
  ram[3438]  = 255;
  ram[3439]  = 255;
  ram[3440]  = 255;
  ram[3441]  = 255;
  ram[3442]  = 255;
  ram[3443]  = 255;
  ram[3444]  = 255;
  ram[3445]  = 255;
  ram[3446]  = 255;
  ram[3447]  = 255;
  ram[3448]  = 255;
  ram[3449]  = 255;
  ram[3450]  = 255;
  ram[3451]  = 255;
  ram[3452]  = 255;
  ram[3453]  = 255;
  ram[3454]  = 255;
  ram[3455]  = 255;
  ram[3456]  = 255;
  ram[3457]  = 255;
  ram[3458]  = 255;
  ram[3459]  = 255;
  ram[3460]  = 255;
  ram[3461]  = 254;
  ram[3462]  = 255;
  ram[3463]  = 110;
  ram[3464]  = 0;
  ram[3465]  = 255;
  ram[3466]  = 255;
  ram[3467]  = 255;
  ram[3468]  = 255;
  ram[3469]  = 255;
  ram[3470]  = 255;
  ram[3471]  = 255;
  ram[3472]  = 255;
  ram[3473]  = 255;
  ram[3474]  = 255;
  ram[3475]  = 255;
  ram[3476]  = 255;
  ram[3477]  = 255;
  ram[3478]  = 255;
  ram[3479]  = 255;
  ram[3480]  = 255;
  ram[3481]  = 255;
  ram[3482]  = 255;
  ram[3483]  = 255;
  ram[3484]  = 255;
  ram[3485]  = 134;
  ram[3486]  = 0;
  ram[3487]  = 246;
  ram[3488]  = 255;
  ram[3489]  = 255;
  ram[3490]  = 255;
  ram[3491]  = 255;
  ram[3492]  = 255;
  ram[3493]  = 255;
  ram[3494]  = 255;
  ram[3495]  = 255;
  ram[3496]  = 255;
  ram[3497]  = 255;
  ram[3498]  = 255;
  ram[3499]  = 255;
  ram[3500]  = 255;
  ram[3501]  = 255;
  ram[3502]  = 255;
  ram[3503]  = 255;
  ram[3504]  = 255;
  ram[3505]  = 255;
  ram[3506]  = 255;
  ram[3507]  = 255;
  ram[3508]  = 255;
  ram[3509]  = 255;
  ram[3510]  = 255;
  ram[3511]  = 255;
  ram[3512]  = 255;
  ram[3513]  = 255;
  ram[3514]  = 255;
  ram[3515]  = 255;
  ram[3516]  = 255;
  ram[3517]  = 255;
  ram[3518]  = 255;
  ram[3519]  = 255;
  ram[3520]  = 255;
  ram[3521]  = 255;
  ram[3522]  = 255;
  ram[3523]  = 255;
  ram[3524]  = 255;
  ram[3525]  = 255;
  ram[3526]  = 255;
  ram[3527]  = 255;
  ram[3528]  = 255;
  ram[3529]  = 255;
  ram[3530]  = 255;
  ram[3531]  = 255;
  ram[3532]  = 255;
  ram[3533]  = 255;
  ram[3534]  = 255;
  ram[3535]  = 255;
  ram[3536]  = 255;
  ram[3537]  = 255;
  ram[3538]  = 255;
  ram[3539]  = 255;
  ram[3540]  = 255;
  ram[3541]  = 255;
  ram[3542]  = 255;
  ram[3543]  = 255;
  ram[3544]  = 255;
  ram[3545]  = 255;
  ram[3546]  = 255;
  ram[3547]  = 255;
  ram[3548]  = 255;
  ram[3549]  = 255;
  ram[3550]  = 255;
  ram[3551]  = 255;
  ram[3552]  = 255;
  ram[3553]  = 255;
  ram[3554]  = 255;
  ram[3555]  = 255;
  ram[3556]  = 255;
  ram[3557]  = 255;
  ram[3558]  = 255;
  ram[3559]  = 255;
  ram[3560]  = 255;
  ram[3561]  = 255;
  ram[3562]  = 255;
  ram[3563]  = 255;
  ram[3564]  = 255;
  ram[3565]  = 255;
  ram[3566]  = 255;
  ram[3567]  = 255;
  ram[3568]  = 255;
  ram[3569]  = 255;
  ram[3570]  = 255;
  ram[3571]  = 255;
  ram[3572]  = 255;
  ram[3573]  = 255;
  ram[3574]  = 255;
  ram[3575]  = 255;
  ram[3576]  = 255;
  ram[3577]  = 255;
  ram[3578]  = 255;
  ram[3579]  = 255;
  ram[3580]  = 255;
  ram[3581]  = 255;
  ram[3582]  = 255;
  ram[3583]  = 255;
  ram[3584]  = 255;
  ram[3585]  = 255;
  ram[3586]  = 255;
  ram[3587]  = 255;
  ram[3588]  = 255;
  ram[3589]  = 255;
  ram[3590]  = 255;
  ram[3591]  = 255;
  ram[3592]  = 255;
  ram[3593]  = 255;
  ram[3594]  = 255;
  ram[3595]  = 255;
  ram[3596]  = 236;
  ram[3597]  = 211;
  ram[3598]  = 243;
  ram[3599]  = 255;
  ram[3600]  = 253;
  ram[3601]  = 235;
  ram[3602]  = 209;
  ram[3603]  = 242;
  ram[3604]  = 255;
  ram[3605]  = 254;
  ram[3606]  = 252;
  ram[3607]  = 255;
  ram[3608]  = 255;
  ram[3609]  = 255;
  ram[3610]  = 255;
  ram[3611]  = 255;
  ram[3612]  = 255;
  ram[3613]  = 255;
  ram[3614]  = 255;
  ram[3615]  = 255;
  ram[3616]  = 167;
  ram[3617]  = 0;
  ram[3618]  = 0;
  ram[3619]  = 0;
  ram[3620]  = 0;
  ram[3621]  = 0;
  ram[3622]  = 151;
  ram[3623]  = 255;
  ram[3624]  = 254;
  ram[3625]  = 255;
  ram[3626]  = 255;
  ram[3627]  = 254;
  ram[3628]  = 254;
  ram[3629]  = 255;
  ram[3630]  = 254;
  ram[3631]  = 254;
  ram[3632]  = 254;
  ram[3633]  = 255;
  ram[3634]  = 254;
  ram[3635]  = 254;
  ram[3636]  = 254;
  ram[3637]  = 255;
  ram[3638]  = 255;
  ram[3639]  = 255;
  ram[3640]  = 255;
  ram[3641]  = 254;
  ram[3642]  = 253;
  ram[3643]  = 254;
  ram[3644]  = 255;
  ram[3645]  = 255;
  ram[3646]  = 255;
  ram[3647]  = 254;
  ram[3648]  = 254;
  ram[3649]  = 254;
  ram[3650]  = 255;
  ram[3651]  = 254;
  ram[3652]  = 255;
  ram[3653]  = 255;
  ram[3654]  = 255;
  ram[3655]  = 255;
  ram[3656]  = 255;
  ram[3657]  = 255;
  ram[3658]  = 255;
  ram[3659]  = 221;
  ram[3660]  = 255;
  ram[3661]  = 254;
  ram[3662]  = 255;
  ram[3663]  = 118;
  ram[3664]  = 0;
  ram[3665]  = 255;
  ram[3666]  = 255;
  ram[3667]  = 254;
  ram[3668]  = 253;
  ram[3669]  = 254;
  ram[3670]  = 255;
  ram[3671]  = 255;
  ram[3672]  = 255;
  ram[3673]  = 255;
  ram[3674]  = 254;
  ram[3675]  = 254;
  ram[3676]  = 254;
  ram[3677]  = 254;
  ram[3678]  = 254;
  ram[3679]  = 255;
  ram[3680]  = 255;
  ram[3681]  = 255;
  ram[3682]  = 255;
  ram[3683]  = 255;
  ram[3684]  = 255;
  ram[3685]  = 144;
  ram[3686]  = 0;
  ram[3687]  = 250;
  ram[3688]  = 255;
  ram[3689]  = 255;
  ram[3690]  = 254;
  ram[3691]  = 254;
  ram[3692]  = 255;
  ram[3693]  = 255;
  ram[3694]  = 255;
  ram[3695]  = 255;
  ram[3696]  = 255;
  ram[3697]  = 255;
  ram[3698]  = 255;
  ram[3699]  = 255;
  ram[3700]  = 255;
  ram[3701]  = 255;
  ram[3702]  = 255;
  ram[3703]  = 255;
  ram[3704]  = 255;
  ram[3705]  = 229;
  ram[3706]  = 250;
  ram[3707]  = 255;
  ram[3708]  = 255;
  ram[3709]  = 255;
  ram[3710]  = 255;
  ram[3711]  = 222;
  ram[3712]  = 255;
  ram[3713]  = 254;
  ram[3714]  = 255;
  ram[3715]  = 255;
  ram[3716]  = 254;
  ram[3717]  = 254;
  ram[3718]  = 254;
  ram[3719]  = 254;
  ram[3720]  = 254;
  ram[3721]  = 255;
  ram[3722]  = 255;
  ram[3723]  = 255;
  ram[3724]  = 255;
  ram[3725]  = 255;
  ram[3726]  = 254;
  ram[3727]  = 255;
  ram[3728]  = 254;
  ram[3729]  = 254;
  ram[3730]  = 254;
  ram[3731]  = 254;
  ram[3732]  = 255;
  ram[3733]  = 255;
  ram[3734]  = 255;
  ram[3735]  = 255;
  ram[3736]  = 255;
  ram[3737]  = 255;
  ram[3738]  = 255;
  ram[3739]  = 245;
  ram[3740]  = 235;
  ram[3741]  = 255;
  ram[3742]  = 255;
  ram[3743]  = 255;
  ram[3744]  = 255;
  ram[3745]  = 255;
  ram[3746]  = 255;
  ram[3747]  = 254;
  ram[3748]  = 254;
  ram[3749]  = 255;
  ram[3750]  = 255;
  ram[3751]  = 255;
  ram[3752]  = 255;
  ram[3753]  = 255;
  ram[3754]  = 255;
  ram[3755]  = 255;
  ram[3756]  = 255;
  ram[3757]  = 255;
  ram[3758]  = 255;
  ram[3759]  = 254;
  ram[3760]  = 254;
  ram[3761]  = 254;
  ram[3762]  = 255;
  ram[3763]  = 254;
  ram[3764]  = 255;
  ram[3765]  = 255;
  ram[3766]  = 222;
  ram[3767]  = 255;
  ram[3768]  = 254;
  ram[3769]  = 255;
  ram[3770]  = 255;
  ram[3771]  = 254;
  ram[3772]  = 254;
  ram[3773]  = 255;
  ram[3774]  = 254;
  ram[3775]  = 255;
  ram[3776]  = 255;
  ram[3777]  = 255;
  ram[3778]  = 255;
  ram[3779]  = 255;
  ram[3780]  = 255;
  ram[3781]  = 254;
  ram[3782]  = 254;
  ram[3783]  = 253;
  ram[3784]  = 255;
  ram[3785]  = 237;
  ram[3786]  = 243;
  ram[3787]  = 255;
  ram[3788]  = 254;
  ram[3789]  = 255;
  ram[3790]  = 255;
  ram[3791]  = 255;
  ram[3792]  = 255;
  ram[3793]  = 255;
  ram[3794]  = 255;
  ram[3795]  = 255;
  ram[3796]  = 235;
  ram[3797]  = 212;
  ram[3798]  = 243;
  ram[3799]  = 255;
  ram[3800]  = 253;
  ram[3801]  = 235;
  ram[3802]  = 209;
  ram[3803]  = 242;
  ram[3804]  = 255;
  ram[3805]  = 254;
  ram[3806]  = 252;
  ram[3807]  = 255;
  ram[3808]  = 255;
  ram[3809]  = 255;
  ram[3810]  = 255;
  ram[3811]  = 255;
  ram[3812]  = 255;
  ram[3813]  = 255;
  ram[3814]  = 255;
  ram[3815]  = 255;
  ram[3816]  = 171;
  ram[3817]  = 0;
  ram[3818]  = 159;
  ram[3819]  = 176;
  ram[3820]  = 158;
  ram[3821]  = 1;
  ram[3822]  = 0;
  ram[3823]  = 219;
  ram[3824]  = 255;
  ram[3825]  = 255;
  ram[3826]  = 255;
  ram[3827]  = 253;
  ram[3828]  = 253;
  ram[3829]  = 254;
  ram[3830]  = 254;
  ram[3831]  = 253;
  ram[3832]  = 253;
  ram[3833]  = 252;
  ram[3834]  = 252;
  ram[3835]  = 253;
  ram[3836]  = 254;
  ram[3837]  = 255;
  ram[3838]  = 255;
  ram[3839]  = 255;
  ram[3840]  = 254;
  ram[3841]  = 254;
  ram[3842]  = 254;
  ram[3843]  = 253;
  ram[3844]  = 254;
  ram[3845]  = 255;
  ram[3846]  = 255;
  ram[3847]  = 253;
  ram[3848]  = 253;
  ram[3849]  = 253;
  ram[3850]  = 252;
  ram[3851]  = 254;
  ram[3852]  = 255;
  ram[3853]  = 255;
  ram[3854]  = 255;
  ram[3855]  = 255;
  ram[3856]  = 254;
  ram[3857]  = 255;
  ram[3858]  = 128;
  ram[3859]  = 11;
  ram[3860]  = 255;
  ram[3861]  = 253;
  ram[3862]  = 255;
  ram[3863]  = 117;
  ram[3864]  = 0;
  ram[3865]  = 255;
  ram[3866]  = 255;
  ram[3867]  = 253;
  ram[3868]  = 253;
  ram[3869]  = 254;
  ram[3870]  = 255;
  ram[3871]  = 255;
  ram[3872]  = 255;
  ram[3873]  = 255;
  ram[3874]  = 253;
  ram[3875]  = 253;
  ram[3876]  = 253;
  ram[3877]  = 254;
  ram[3878]  = 253;
  ram[3879]  = 255;
  ram[3880]  = 255;
  ram[3881]  = 255;
  ram[3882]  = 255;
  ram[3883]  = 255;
  ram[3884]  = 255;
  ram[3885]  = 141;
  ram[3886]  = 0;
  ram[3887]  = 250;
  ram[3888]  = 255;
  ram[3889]  = 253;
  ram[3890]  = 252;
  ram[3891]  = 253;
  ram[3892]  = 255;
  ram[3893]  = 255;
  ram[3894]  = 255;
  ram[3895]  = 255;
  ram[3896]  = 255;
  ram[3897]  = 255;
  ram[3898]  = 255;
  ram[3899]  = 255;
  ram[3900]  = 255;
  ram[3901]  = 255;
  ram[3902]  = 255;
  ram[3903]  = 255;
  ram[3904]  = 204;
  ram[3905]  = 0;
  ram[3906]  = 240;
  ram[3907]  = 255;
  ram[3908]  = 255;
  ram[3909]  = 255;
  ram[3910]  = 93;
  ram[3911]  = 43;
  ram[3912]  = 255;
  ram[3913]  = 251;
  ram[3914]  = 255;
  ram[3915]  = 255;
  ram[3916]  = 254;
  ram[3917]  = 253;
  ram[3918]  = 253;
  ram[3919]  = 253;
  ram[3920]  = 254;
  ram[3921]  = 255;
  ram[3922]  = 255;
  ram[3923]  = 255;
  ram[3924]  = 255;
  ram[3925]  = 255;
  ram[3926]  = 254;
  ram[3927]  = 252;
  ram[3928]  = 253;
  ram[3929]  = 253;
  ram[3930]  = 253;
  ram[3931]  = 254;
  ram[3932]  = 255;
  ram[3933]  = 255;
  ram[3934]  = 255;
  ram[3935]  = 255;
  ram[3936]  = 255;
  ram[3937]  = 255;
  ram[3938]  = 247;
  ram[3939]  = 12;
  ram[3940]  = 159;
  ram[3941]  = 255;
  ram[3942]  = 255;
  ram[3943]  = 255;
  ram[3944]  = 255;
  ram[3945]  = 255;
  ram[3946]  = 253;
  ram[3947]  = 252;
  ram[3948]  = 254;
  ram[3949]  = 255;
  ram[3950]  = 255;
  ram[3951]  = 255;
  ram[3952]  = 255;
  ram[3953]  = 255;
  ram[3954]  = 255;
  ram[3955]  = 255;
  ram[3956]  = 255;
  ram[3957]  = 255;
  ram[3958]  = 254;
  ram[3959]  = 253;
  ram[3960]  = 255;
  ram[3961]  = 253;
  ram[3962]  = 253;
  ram[3963]  = 253;
  ram[3964]  = 255;
  ram[3965]  = 95;
  ram[3966]  = 44;
  ram[3967]  = 255;
  ram[3968]  = 254;
  ram[3969]  = 255;
  ram[3970]  = 255;
  ram[3971]  = 253;
  ram[3972]  = 253;
  ram[3973]  = 253;
  ram[3974]  = 253;
  ram[3975]  = 255;
  ram[3976]  = 255;
  ram[3977]  = 255;
  ram[3978]  = 255;
  ram[3979]  = 255;
  ram[3980]  = 255;
  ram[3981]  = 252;
  ram[3982]  = 252;
  ram[3983]  = 255;
  ram[3984]  = 224;
  ram[3985]  = 0;
  ram[3986]  = 202;
  ram[3987]  = 255;
  ram[3988]  = 253;
  ram[3989]  = 255;
  ram[3990]  = 255;
  ram[3991]  = 255;
  ram[3992]  = 255;
  ram[3993]  = 255;
  ram[3994]  = 255;
  ram[3995]  = 255;
  ram[3996]  = 235;
  ram[3997]  = 212;
  ram[3998]  = 243;
  ram[3999]  = 255;
  ram[4000]  = 253;
  ram[4001]  = 235;
  ram[4002]  = 209;
  ram[4003]  = 242;
  ram[4004]  = 255;
  ram[4005]  = 254;
  ram[4006]  = 252;
  ram[4007]  = 255;
  ram[4008]  = 255;
  ram[4009]  = 255;
  ram[4010]  = 255;
  ram[4011]  = 255;
  ram[4012]  = 255;
  ram[4013]  = 255;
  ram[4014]  = 255;
  ram[4015]  = 255;
  ram[4016]  = 170;
  ram[4017]  = 0;
  ram[4018]  = 238;
  ram[4019]  = 255;
  ram[4020]  = 255;
  ram[4021]  = 237;
  ram[4022]  = 0;
  ram[4023]  = 114;
  ram[4024]  = 255;
  ram[4025]  = 255;
  ram[4026]  = 255;
  ram[4027]  = 255;
  ram[4028]  = 255;
  ram[4029]  = 255;
  ram[4030]  = 252;
  ram[4031]  = 254;
  ram[4032]  = 254;
  ram[4033]  = 255;
  ram[4034]  = 255;
  ram[4035]  = 255;
  ram[4036]  = 255;
  ram[4037]  = 255;
  ram[4038]  = 255;
  ram[4039]  = 254;
  ram[4040]  = 255;
  ram[4041]  = 255;
  ram[4042]  = 255;
  ram[4043]  = 255;
  ram[4044]  = 255;
  ram[4045]  = 255;
  ram[4046]  = 255;
  ram[4047]  = 255;
  ram[4048]  = 255;
  ram[4049]  = 255;
  ram[4050]  = 255;
  ram[4051]  = 254;
  ram[4052]  = 255;
  ram[4053]  = 255;
  ram[4054]  = 255;
  ram[4055]  = 255;
  ram[4056]  = 254;
  ram[4057]  = 255;
  ram[4058]  = 83;
  ram[4059]  = 8;
  ram[4060]  = 255;
  ram[4061]  = 255;
  ram[4062]  = 255;
  ram[4063]  = 117;
  ram[4064]  = 0;
  ram[4065]  = 255;
  ram[4066]  = 255;
  ram[4067]  = 255;
  ram[4068]  = 255;
  ram[4069]  = 255;
  ram[4070]  = 255;
  ram[4071]  = 255;
  ram[4072]  = 255;
  ram[4073]  = 254;
  ram[4074]  = 255;
  ram[4075]  = 255;
  ram[4076]  = 255;
  ram[4077]  = 255;
  ram[4078]  = 253;
  ram[4079]  = 255;
  ram[4080]  = 255;
  ram[4081]  = 255;
  ram[4082]  = 255;
  ram[4083]  = 255;
  ram[4084]  = 255;
  ram[4085]  = 141;
  ram[4086]  = 0;
  ram[4087]  = 250;
  ram[4088]  = 255;
  ram[4089]  = 255;
  ram[4090]  = 255;
  ram[4091]  = 255;
  ram[4092]  = 255;
  ram[4093]  = 255;
  ram[4094]  = 255;
  ram[4095]  = 255;
  ram[4096]  = 255;
  ram[4097]  = 255;
  ram[4098]  = 255;
  ram[4099]  = 255;
  ram[4100]  = 255;
  ram[4101]  = 255;
  ram[4102]  = 255;
  ram[4103]  = 255;
  ram[4104]  = 181;
  ram[4105]  = 0;
  ram[4106]  = 251;
  ram[4107]  = 255;
  ram[4108]  = 255;
  ram[4109]  = 255;
  ram[4110]  = 42;
  ram[4111]  = 49;
  ram[4112]  = 255;
  ram[4113]  = 254;
  ram[4114]  = 255;
  ram[4115]  = 255;
  ram[4116]  = 255;
  ram[4117]  = 255;
  ram[4118]  = 255;
  ram[4119]  = 255;
  ram[4120]  = 255;
  ram[4121]  = 255;
  ram[4122]  = 255;
  ram[4123]  = 255;
  ram[4124]  = 255;
  ram[4125]  = 255;
  ram[4126]  = 255;
  ram[4127]  = 255;
  ram[4128]  = 255;
  ram[4129]  = 255;
  ram[4130]  = 255;
  ram[4131]  = 255;
  ram[4132]  = 255;
  ram[4133]  = 255;
  ram[4134]  = 255;
  ram[4135]  = 255;
  ram[4136]  = 255;
  ram[4137]  = 255;
  ram[4138]  = 246;
  ram[4139]  = 0;
  ram[4140]  = 170;
  ram[4141]  = 255;
  ram[4142]  = 255;
  ram[4143]  = 255;
  ram[4144]  = 255;
  ram[4145]  = 255;
  ram[4146]  = 255;
  ram[4147]  = 255;
  ram[4148]  = 255;
  ram[4149]  = 255;
  ram[4150]  = 254;
  ram[4151]  = 255;
  ram[4152]  = 255;
  ram[4153]  = 255;
  ram[4154]  = 255;
  ram[4155]  = 255;
  ram[4156]  = 255;
  ram[4157]  = 255;
  ram[4158]  = 255;
  ram[4159]  = 255;
  ram[4160]  = 255;
  ram[4161]  = 255;
  ram[4162]  = 255;
  ram[4163]  = 254;
  ram[4164]  = 255;
  ram[4165]  = 41;
  ram[4166]  = 50;
  ram[4167]  = 255;
  ram[4168]  = 255;
  ram[4169]  = 255;
  ram[4170]  = 255;
  ram[4171]  = 255;
  ram[4172]  = 255;
  ram[4173]  = 255;
  ram[4174]  = 255;
  ram[4175]  = 254;
  ram[4176]  = 254;
  ram[4177]  = 255;
  ram[4178]  = 255;
  ram[4179]  = 255;
  ram[4180]  = 255;
  ram[4181]  = 255;
  ram[4182]  = 255;
  ram[4183]  = 255;
  ram[4184]  = 209;
  ram[4185]  = 0;
  ram[4186]  = 215;
  ram[4187]  = 255;
  ram[4188]  = 255;
  ram[4189]  = 255;
  ram[4190]  = 255;
  ram[4191]  = 255;
  ram[4192]  = 255;
  ram[4193]  = 255;
  ram[4194]  = 255;
  ram[4195]  = 255;
  ram[4196]  = 236;
  ram[4197]  = 211;
  ram[4198]  = 243;
  ram[4199]  = 255;
  ram[4200]  = 253;
  ram[4201]  = 235;
  ram[4202]  = 209;
  ram[4203]  = 242;
  ram[4204]  = 255;
  ram[4205]  = 254;
  ram[4206]  = 252;
  ram[4207]  = 255;
  ram[4208]  = 255;
  ram[4209]  = 255;
  ram[4210]  = 255;
  ram[4211]  = 255;
  ram[4212]  = 255;
  ram[4213]  = 255;
  ram[4214]  = 255;
  ram[4215]  = 255;
  ram[4216]  = 170;
  ram[4217]  = 0;
  ram[4218]  = 229;
  ram[4219]  = 255;
  ram[4220]  = 253;
  ram[4221]  = 255;
  ram[4222]  = 19;
  ram[4223]  = 63;
  ram[4224]  = 255;
  ram[4225]  = 243;
  ram[4226]  = 219;
  ram[4227]  = 255;
  ram[4228]  = 206;
  ram[4229]  = 185;
  ram[4230]  = 255;
  ram[4231]  = 255;
  ram[4232]  = 255;
  ram[4233]  = 203;
  ram[4234]  = 152;
  ram[4235]  = 205;
  ram[4236]  = 255;
  ram[4237]  = 255;
  ram[4238]  = 254;
  ram[4239]  = 255;
  ram[4240]  = 253;
  ram[4241]  = 190;
  ram[4242]  = 153;
  ram[4243]  = 199;
  ram[4244]  = 253;
  ram[4245]  = 255;
  ram[4246]  = 255;
  ram[4247]  = 251;
  ram[4248]  = 183;
  ram[4249]  = 152;
  ram[4250]  = 203;
  ram[4251]  = 255;
  ram[4252]  = 255;
  ram[4253]  = 255;
  ram[4254]  = 255;
  ram[4255]  = 255;
  ram[4256]  = 255;
  ram[4257]  = 240;
  ram[4258]  = 77;
  ram[4259]  = 10;
  ram[4260]  = 245;
  ram[4261]  = 228;
  ram[4262]  = 255;
  ram[4263]  = 117;
  ram[4264]  = 0;
  ram[4265]  = 255;
  ram[4266]  = 217;
  ram[4267]  = 150;
  ram[4268]  = 199;
  ram[4269]  = 255;
  ram[4270]  = 255;
  ram[4271]  = 253;
  ram[4272]  = 254;
  ram[4273]  = 255;
  ram[4274]  = 235;
  ram[4275]  = 166;
  ram[4276]  = 168;
  ram[4277]  = 243;
  ram[4278]  = 255;
  ram[4279]  = 255;
  ram[4280]  = 255;
  ram[4281]  = 255;
  ram[4282]  = 255;
  ram[4283]  = 255;
  ram[4284]  = 255;
  ram[4285]  = 141;
  ram[4286]  = 0;
  ram[4287]  = 255;
  ram[4288]  = 233;
  ram[4289]  = 153;
  ram[4290]  = 185;
  ram[4291]  = 255;
  ram[4292]  = 255;
  ram[4293]  = 255;
  ram[4294]  = 255;
  ram[4295]  = 217;
  ram[4296]  = 245;
  ram[4297]  = 255;
  ram[4298]  = 255;
  ram[4299]  = 255;
  ram[4300]  = 229;
  ram[4301]  = 229;
  ram[4302]  = 255;
  ram[4303]  = 241;
  ram[4304]  = 157;
  ram[4305]  = 0;
  ram[4306]  = 216;
  ram[4307]  = 228;
  ram[4308]  = 253;
  ram[4309]  = 241;
  ram[4310]  = 44;
  ram[4311]  = 43;
  ram[4312]  = 241;
  ram[4313]  = 233;
  ram[4314]  = 255;
  ram[4315]  = 255;
  ram[4316]  = 255;
  ram[4317]  = 225;
  ram[4318]  = 159;
  ram[4319]  = 168;
  ram[4320]  = 233;
  ram[4321]  = 255;
  ram[4322]  = 255;
  ram[4323]  = 255;
  ram[4324]  = 252;
  ram[4325]  = 217;
  ram[4326]  = 255;
  ram[4327]  = 244;
  ram[4328]  = 161;
  ram[4329]  = 178;
  ram[4330]  = 251;
  ram[4331]  = 255;
  ram[4332]  = 254;
  ram[4333]  = 254;
  ram[4334]  = 255;
  ram[4335]  = 255;
  ram[4336]  = 255;
  ram[4337]  = 247;
  ram[4338]  = 209;
  ram[4339]  = 0;
  ram[4340]  = 146;
  ram[4341]  = 231;
  ram[4342]  = 245;
  ram[4343]  = 255;
  ram[4344]  = 255;
  ram[4345]  = 255;
  ram[4346]  = 196;
  ram[4347]  = 151;
  ram[4348]  = 183;
  ram[4349]  = 254;
  ram[4350]  = 255;
  ram[4351]  = 254;
  ram[4352]  = 254;
  ram[4353]  = 255;
  ram[4354]  = 255;
  ram[4355]  = 255;
  ram[4356]  = 254;
  ram[4357]  = 255;
  ram[4358]  = 255;
  ram[4359]  = 205;
  ram[4360]  = 153;
  ram[4361]  = 183;
  ram[4362]  = 246;
  ram[4363]  = 255;
  ram[4364]  = 241;
  ram[4365]  = 44;
  ram[4366]  = 44;
  ram[4367]  = 241;
  ram[4368]  = 233;
  ram[4369]  = 255;
  ram[4370]  = 255;
  ram[4371]  = 241;
  ram[4372]  = 178;
  ram[4373]  = 155;
  ram[4374]  = 214;
  ram[4375]  = 255;
  ram[4376]  = 255;
  ram[4377]  = 255;
  ram[4378]  = 245;
  ram[4379]  = 219;
  ram[4380]  = 255;
  ram[4381]  = 209;
  ram[4382]  = 183;
  ram[4383]  = 250;
  ram[4384]  = 180;
  ram[4385]  = 0;
  ram[4386]  = 183;
  ram[4387]  = 227;
  ram[4388]  = 252;
  ram[4389]  = 255;
  ram[4390]  = 255;
  ram[4391]  = 255;
  ram[4392]  = 255;
  ram[4393]  = 255;
  ram[4394]  = 255;
  ram[4395]  = 255;
  ram[4396]  = 236;
  ram[4397]  = 211;
  ram[4398]  = 243;
  ram[4399]  = 255;
  ram[4400]  = 253;
  ram[4401]  = 235;
  ram[4402]  = 209;
  ram[4403]  = 242;
  ram[4404]  = 255;
  ram[4405]  = 254;
  ram[4406]  = 252;
  ram[4407]  = 255;
  ram[4408]  = 255;
  ram[4409]  = 255;
  ram[4410]  = 255;
  ram[4411]  = 255;
  ram[4412]  = 255;
  ram[4413]  = 255;
  ram[4414]  = 255;
  ram[4415]  = 255;
  ram[4416]  = 170;
  ram[4417]  = 0;
  ram[4418]  = 231;
  ram[4419]  = 255;
  ram[4420]  = 253;
  ram[4421]  = 255;
  ram[4422]  = 29;
  ram[4423]  = 65;
  ram[4424]  = 255;
  ram[4425]  = 151;
  ram[4426]  = 0;
  ram[4427]  = 181;
  ram[4428]  = 0;
  ram[4429]  = 0;
  ram[4430]  = 255;
  ram[4431]  = 255;
  ram[4432]  = 106;
  ram[4433]  = 0;
  ram[4434]  = 0;
  ram[4435]  = 0;
  ram[4436]  = 123;
  ram[4437]  = 255;
  ram[4438]  = 255;
  ram[4439]  = 255;
  ram[4440]  = 53;
  ram[4441]  = 0;
  ram[4442]  = 0;
  ram[4443]  = 0;
  ram[4444]  = 190;
  ram[4445]  = 255;
  ram[4446]  = 253;
  ram[4447]  = 35;
  ram[4448]  = 0;
  ram[4449]  = 0;
  ram[4450]  = 0;
  ram[4451]  = 226;
  ram[4452]  = 255;
  ram[4453]  = 255;
  ram[4454]  = 255;
  ram[4455]  = 255;
  ram[4456]  = 249;
  ram[4457]  = 0;
  ram[4458]  = 0;
  ram[4459]  = 0;
  ram[4460]  = 0;
  ram[4461]  = 29;
  ram[4462]  = 255;
  ram[4463]  = 118;
  ram[4464]  = 15;
  ram[4465]  = 187;
  ram[4466]  = 0;
  ram[4467]  = 0;
  ram[4468]  = 0;
  ram[4469]  = 154;
  ram[4470]  = 255;
  ram[4471]  = 251;
  ram[4472]  = 255;
  ram[4473]  = 216;
  ram[4474]  = 5;
  ram[4475]  = 0;
  ram[4476]  = 0;
  ram[4477]  = 21;
  ram[4478]  = 240;
  ram[4479]  = 255;
  ram[4480]  = 255;
  ram[4481]  = 255;
  ram[4482]  = 255;
  ram[4483]  = 255;
  ram[4484]  = 255;
  ram[4485]  = 141;
  ram[4486]  = 3;
  ram[4487]  = 195;
  ram[4488]  = 0;
  ram[4489]  = 0;
  ram[4490]  = 0;
  ram[4491]  = 76;
  ram[4492]  = 255;
  ram[4493]  = 255;
  ram[4494]  = 245;
  ram[4495]  = 0;
  ram[4496]  = 169;
  ram[4497]  = 255;
  ram[4498]  = 255;
  ram[4499]  = 255;
  ram[4500]  = 57;
  ram[4501]  = 40;
  ram[4502]  = 255;
  ram[4503]  = 66;
  ram[4504]  = 0;
  ram[4505]  = 0;
  ram[4506]  = 0;
  ram[4507]  = 0;
  ram[4508]  = 206;
  ram[4509]  = 0;
  ram[4510]  = 0;
  ram[4511]  = 0;
  ram[4512]  = 0;
  ram[4513]  = 61;
  ram[4514]  = 255;
  ram[4515]  = 255;
  ram[4516]  = 144;
  ram[4517]  = 0;
  ram[4518]  = 0;
  ram[4519]  = 0;
  ram[4520]  = 0;
  ram[4521]  = 188;
  ram[4522]  = 255;
  ram[4523]  = 255;
  ram[4524]  = 222;
  ram[4525]  = 0;
  ram[4526]  = 189;
  ram[4527]  = 19;
  ram[4528]  = 0;
  ram[4529]  = 0;
  ram[4530]  = 63;
  ram[4531]  = 255;
  ram[4532]  = 254;
  ram[4533]  = 252;
  ram[4534]  = 255;
  ram[4535]  = 255;
  ram[4536]  = 255;
  ram[4537]  = 146;
  ram[4538]  = 0;
  ram[4539]  = 0;
  ram[4540]  = 0;
  ram[4541]  = 0;
  ram[4542]  = 158;
  ram[4543]  = 255;
  ram[4544]  = 255;
  ram[4545]  = 62;
  ram[4546]  = 0;
  ram[4547]  = 0;
  ram[4548]  = 0;
  ram[4549]  = 41;
  ram[4550]  = 247;
  ram[4551]  = 255;
  ram[4552]  = 254;
  ram[4553]  = 254;
  ram[4554]  = 255;
  ram[4555]  = 255;
  ram[4556]  = 248;
  ram[4557]  = 255;
  ram[4558]  = 104;
  ram[4559]  = 0;
  ram[4560]  = 0;
  ram[4561]  = 0;
  ram[4562]  = 118;
  ram[4563]  = 245;
  ram[4564]  = 0;
  ram[4565]  = 0;
  ram[4566]  = 0;
  ram[4567]  = 0;
  ram[4568]  = 62;
  ram[4569]  = 255;
  ram[4570]  = 201;
  ram[4571]  = 1;
  ram[4572]  = 0;
  ram[4573]  = 0;
  ram[4574]  = 0;
  ram[4575]  = 168;
  ram[4576]  = 255;
  ram[4577]  = 255;
  ram[4578]  = 159;
  ram[4579]  = 0;
  ram[4580]  = 180;
  ram[4581]  = 0;
  ram[4582]  = 0;
  ram[4583]  = 121;
  ram[4584]  = 0;
  ram[4585]  = 0;
  ram[4586]  = 0;
  ram[4587]  = 0;
  ram[4588]  = 210;
  ram[4589]  = 255;
  ram[4590]  = 255;
  ram[4591]  = 255;
  ram[4592]  = 255;
  ram[4593]  = 255;
  ram[4594]  = 255;
  ram[4595]  = 255;
  ram[4596]  = 236;
  ram[4597]  = 211;
  ram[4598]  = 243;
  ram[4599]  = 255;
  ram[4600]  = 253;
  ram[4601]  = 235;
  ram[4602]  = 209;
  ram[4603]  = 242;
  ram[4604]  = 255;
  ram[4605]  = 254;
  ram[4606]  = 252;
  ram[4607]  = 255;
  ram[4608]  = 255;
  ram[4609]  = 255;
  ram[4610]  = 255;
  ram[4611]  = 255;
  ram[4612]  = 255;
  ram[4613]  = 255;
  ram[4614]  = 255;
  ram[4615]  = 255;
  ram[4616]  = 170;
  ram[4617]  = 0;
  ram[4618]  = 233;
  ram[4619]  = 255;
  ram[4620]  = 255;
  ram[4621]  = 255;
  ram[4622]  = 0;
  ram[4623]  = 109;
  ram[4624]  = 255;
  ram[4625]  = 153;
  ram[4626]  = 0;
  ram[4627]  = 23;
  ram[4628]  = 133;
  ram[4629]  = 142;
  ram[4630]  = 255;
  ram[4631]  = 157;
  ram[4632]  = 0;
  ram[4633]  = 140;
  ram[4634]  = 245;
  ram[4635]  = 114;
  ram[4636]  = 0;
  ram[4637]  = 215;
  ram[4638]  = 255;
  ram[4639]  = 118;
  ram[4640]  = 0;
  ram[4641]  = 187;
  ram[4642]  = 240;
  ram[4643]  = 146;
  ram[4644]  = 198;
  ram[4645]  = 255;
  ram[4646]  = 88;
  ram[4647]  = 0;
  ram[4648]  = 201;
  ram[4649]  = 239;
  ram[4650]  = 126;
  ram[4651]  = 215;
  ram[4652]  = 255;
  ram[4653]  = 255;
  ram[4654]  = 255;
  ram[4655]  = 255;
  ram[4656]  = 254;
  ram[4657]  = 164;
  ram[4658]  = 52;
  ram[4659]  = 10;
  ram[4660]  = 163;
  ram[4661]  = 168;
  ram[4662]  = 255;
  ram[4663]  = 123;
  ram[4664]  = 0;
  ram[4665]  = 19;
  ram[4666]  = 190;
  ram[4667]  = 222;
  ram[4668]  = 10;
  ram[4669]  = 1;
  ram[4670]  = 253;
  ram[4671]  = 255;
  ram[4672]  = 255;
  ram[4673]  = 1;
  ram[4674]  = 36;
  ram[4675]  = 220;
  ram[4676]  = 215;
  ram[4677]  = 0;
  ram[4678]  = 64;
  ram[4679]  = 255;
  ram[4680]  = 255;
  ram[4681]  = 255;
  ram[4682]  = 255;
  ram[4683]  = 255;
  ram[4684]  = 255;
  ram[4685]  = 143;
  ram[4686]  = 0;
  ram[4687]  = 15;
  ram[4688]  = 155;
  ram[4689]  = 236;
  ram[4690]  = 102;
  ram[4691]  = 0;
  ram[4692]  = 151;
  ram[4693]  = 255;
  ram[4694]  = 247;
  ram[4695]  = 0;
  ram[4696]  = 171;
  ram[4697]  = 255;
  ram[4698]  = 255;
  ram[4699]  = 255;
  ram[4700]  = 60;
  ram[4701]  = 39;
  ram[4702]  = 255;
  ram[4703]  = 189;
  ram[4704]  = 100;
  ram[4705]  = 0;
  ram[4706]  = 147;
  ram[4707]  = 151;
  ram[4708]  = 236;
  ram[4709]  = 160;
  ram[4710]  = 29;
  ram[4711]  = 29;
  ram[4712]  = 160;
  ram[4713]  = 176;
  ram[4714]  = 255;
  ram[4715]  = 196;
  ram[4716]  = 0;
  ram[4717]  = 80;
  ram[4718]  = 222;
  ram[4719]  = 199;
  ram[4720]  = 32;
  ram[4721]  = 0;
  ram[4722]  = 238;
  ram[4723]  = 255;
  ram[4724]  = 226;
  ram[4725]  = 0;
  ram[4726]  = 1;
  ram[4727]  = 131;
  ram[4728]  = 234;
  ram[4729]  = 91;
  ram[4730]  = 0;
  ram[4731]  = 189;
  ram[4732]  = 255;
  ram[4733]  = 253;
  ram[4734]  = 255;
  ram[4735]  = 255;
  ram[4736]  = 255;
  ram[4737]  = 214;
  ram[4738]  = 136;
  ram[4739]  = 0;
  ram[4740]  = 101;
  ram[4741]  = 153;
  ram[4742]  = 214;
  ram[4743]  = 255;
  ram[4744]  = 85;
  ram[4745]  = 0;
  ram[4746]  = 147;
  ram[4747]  = 233;
  ram[4748]  = 163;
  ram[4749]  = 0;
  ram[4750]  = 53;
  ram[4751]  = 255;
  ram[4752]  = 254;
  ram[4753]  = 255;
  ram[4754]  = 255;
  ram[4755]  = 255;
  ram[4756]  = 255;
  ram[4757]  = 189;
  ram[4758]  = 0;
  ram[4759]  = 140;
  ram[4760]  = 244;
  ram[4761]  = 178;
  ram[4762]  = 152;
  ram[4763]  = 255;
  ram[4764]  = 158;
  ram[4765]  = 27;
  ram[4766]  = 31;
  ram[4767]  = 160;
  ram[4768]  = 178;
  ram[4769]  = 255;
  ram[4770]  = 128;
  ram[4771]  = 73;
  ram[4772]  = 216;
  ram[4773]  = 235;
  ram[4774]  = 37;
  ram[4775]  = 0;
  ram[4776]  = 255;
  ram[4777]  = 255;
  ram[4778]  = 162;
  ram[4779]  = 0;
  ram[4780]  = 27;
  ram[4781]  = 128;
  ram[4782]  = 140;
  ram[4783]  = 207;
  ram[4784]  = 116;
  ram[4785]  = 0;
  ram[4786]  = 123;
  ram[4787]  = 146;
  ram[4788]  = 240;
  ram[4789]  = 255;
  ram[4790]  = 255;
  ram[4791]  = 255;
  ram[4792]  = 255;
  ram[4793]  = 255;
  ram[4794]  = 255;
  ram[4795]  = 255;
  ram[4796]  = 236;
  ram[4797]  = 211;
  ram[4798]  = 243;
  ram[4799]  = 255;
  ram[4800]  = 253;
  ram[4801]  = 235;
  ram[4802]  = 209;
  ram[4803]  = 242;
  ram[4804]  = 255;
  ram[4805]  = 254;
  ram[4806]  = 252;
  ram[4807]  = 255;
  ram[4808]  = 255;
  ram[4809]  = 255;
  ram[4810]  = 255;
  ram[4811]  = 255;
  ram[4812]  = 255;
  ram[4813]  = 255;
  ram[4814]  = 255;
  ram[4815]  = 255;
  ram[4816]  = 170;
  ram[4817]  = 0;
  ram[4818]  = 232;
  ram[4819]  = 255;
  ram[4820]  = 254;
  ram[4821]  = 94;
  ram[4822]  = 0;
  ram[4823]  = 201;
  ram[4824]  = 255;
  ram[4825]  = 157;
  ram[4826]  = 0;
  ram[4827]  = 129;
  ram[4828]  = 255;
  ram[4829]  = 255;
  ram[4830]  = 255;
  ram[4831]  = 11;
  ram[4832]  = 85;
  ram[4833]  = 255;
  ram[4834]  = 255;
  ram[4835]  = 255;
  ram[4836]  = 16;
  ram[4837]  = 103;
  ram[4838]  = 255;
  ram[4839]  = 47;
  ram[4840]  = 54;
  ram[4841]  = 255;
  ram[4842]  = 255;
  ram[4843]  = 255;
  ram[4844]  = 255;
  ram[4845]  = 255;
  ram[4846]  = 10;
  ram[4847]  = 75;
  ram[4848]  = 255;
  ram[4849]  = 255;
  ram[4850]  = 255;
  ram[4851]  = 252;
  ram[4852]  = 255;
  ram[4853]  = 255;
  ram[4854]  = 255;
  ram[4855]  = 255;
  ram[4856]  = 255;
  ram[4857]  = 255;
  ram[4858]  = 91;
  ram[4859]  = 11;
  ram[4860]  = 255;
  ram[4861]  = 255;
  ram[4862]  = 255;
  ram[4863]  = 122;
  ram[4864]  = 0;
  ram[4865]  = 179;
  ram[4866]  = 255;
  ram[4867]  = 255;
  ram[4868]  = 171;
  ram[4869]  = 0;
  ram[4870]  = 210;
  ram[4871]  = 255;
  ram[4872]  = 159;
  ram[4873]  = 0;
  ram[4874]  = 232;
  ram[4875]  = 255;
  ram[4876]  = 255;
  ram[4877]  = 170;
  ram[4878]  = 0;
  ram[4879]  = 244;
  ram[4880]  = 255;
  ram[4881]  = 255;
  ram[4882]  = 255;
  ram[4883]  = 255;
  ram[4884]  = 255;
  ram[4885]  = 145;
  ram[4886]  = 0;
  ram[4887]  = 144;
  ram[4888]  = 255;
  ram[4889]  = 255;
  ram[4890]  = 255;
  ram[4891]  = 30;
  ram[4892]  = 32;
  ram[4893]  = 255;
  ram[4894]  = 248;
  ram[4895]  = 0;
  ram[4896]  = 172;
  ram[4897]  = 255;
  ram[4898]  = 255;
  ram[4899]  = 255;
  ram[4900]  = 59;
  ram[4901]  = 40;
  ram[4902]  = 255;
  ram[4903]  = 255;
  ram[4904]  = 188;
  ram[4905]  = 0;
  ram[4906]  = 254;
  ram[4907]  = 255;
  ram[4908]  = 255;
  ram[4909]  = 255;
  ram[4910]  = 52;
  ram[4911]  = 52;
  ram[4912]  = 255;
  ram[4913]  = 255;
  ram[4914]  = 255;
  ram[4915]  = 35;
  ram[4916]  = 32;
  ram[4917]  = 255;
  ram[4918]  = 255;
  ram[4919]  = 255;
  ram[4920]  = 232;
  ram[4921]  = 0;
  ram[4922]  = 131;
  ram[4923]  = 255;
  ram[4924]  = 224;
  ram[4925]  = 0;
  ram[4926]  = 76;
  ram[4927]  = 255;
  ram[4928]  = 255;
  ram[4929]  = 252;
  ram[4930]  = 0;
  ram[4931]  = 107;
  ram[4932]  = 255;
  ram[4933]  = 253;
  ram[4934]  = 255;
  ram[4935]  = 255;
  ram[4936]  = 253;
  ram[4937]  = 255;
  ram[4938]  = 254;
  ram[4939]  = 0;
  ram[4940]  = 177;
  ram[4941]  = 255;
  ram[4942]  = 255;
  ram[4943]  = 238;
  ram[4944]  = 0;
  ram[4945]  = 122;
  ram[4946]  = 255;
  ram[4947]  = 255;
  ram[4948]  = 255;
  ram[4949]  = 145;
  ram[4950]  = 0;
  ram[4951]  = 225;
  ram[4952]  = 255;
  ram[4953]  = 255;
  ram[4954]  = 255;
  ram[4955]  = 255;
  ram[4956]  = 255;
  ram[4957]  = 116;
  ram[4958]  = 0;
  ram[4959]  = 255;
  ram[4960]  = 255;
  ram[4961]  = 255;
  ram[4962]  = 255;
  ram[4963]  = 253;
  ram[4964]  = 255;
  ram[4965]  = 53;
  ram[4966]  = 53;
  ram[4967]  = 255;
  ram[4968]  = 255;
  ram[4969]  = 253;
  ram[4970]  = 233;
  ram[4971]  = 255;
  ram[4972]  = 255;
  ram[4973]  = 255;
  ram[4974]  = 202;
  ram[4975]  = 0;
  ram[4976]  = 219;
  ram[4977]  = 255;
  ram[4978]  = 161;
  ram[4979]  = 0;
  ram[4980]  = 118;
  ram[4981]  = 255;
  ram[4982]  = 255;
  ram[4983]  = 255;
  ram[4984]  = 217;
  ram[4985]  = 0;
  ram[4986]  = 220;
  ram[4987]  = 255;
  ram[4988]  = 255;
  ram[4989]  = 255;
  ram[4990]  = 255;
  ram[4991]  = 255;
  ram[4992]  = 255;
  ram[4993]  = 255;
  ram[4994]  = 255;
  ram[4995]  = 255;
  ram[4996]  = 235;
  ram[4997]  = 211;
  ram[4998]  = 243;
  ram[4999]  = 255;
  ram[5000]  = 253;
  ram[5001]  = 235;
  ram[5002]  = 209;
  ram[5003]  = 242;
  ram[5004]  = 255;
  ram[5005]  = 254;
  ram[5006]  = 252;
  ram[5007]  = 255;
  ram[5008]  = 255;
  ram[5009]  = 255;
  ram[5010]  = 255;
  ram[5011]  = 255;
  ram[5012]  = 255;
  ram[5013]  = 255;
  ram[5014]  = 255;
  ram[5015]  = 255;
  ram[5016]  = 171;
  ram[5017]  = 0;
  ram[5018]  = 48;
  ram[5019]  = 50;
  ram[5020]  = 22;
  ram[5021]  = 0;
  ram[5022]  = 88;
  ram[5023]  = 255;
  ram[5024]  = 255;
  ram[5025]  = 155;
  ram[5026]  = 0;
  ram[5027]  = 220;
  ram[5028]  = 255;
  ram[5029]  = 255;
  ram[5030]  = 232;
  ram[5031]  = 0;
  ram[5032]  = 200;
  ram[5033]  = 255;
  ram[5034]  = 255;
  ram[5035]  = 255;
  ram[5036]  = 73;
  ram[5037]  = 42;
  ram[5038]  = 255;
  ram[5039]  = 71;
  ram[5040]  = 0;
  ram[5041]  = 232;
  ram[5042]  = 255;
  ram[5043]  = 255;
  ram[5044]  = 251;
  ram[5045]  = 255;
  ram[5046]  = 37;
  ram[5047]  = 13;
  ram[5048]  = 245;
  ram[5049]  = 255;
  ram[5050]  = 254;
  ram[5051]  = 252;
  ram[5052]  = 254;
  ram[5053]  = 254;
  ram[5054]  = 255;
  ram[5055]  = 255;
  ram[5056]  = 254;
  ram[5057]  = 255;
  ram[5058]  = 86;
  ram[5059]  = 8;
  ram[5060]  = 255;
  ram[5061]  = 255;
  ram[5062]  = 255;
  ram[5063]  = 119;
  ram[5064]  = 0;
  ram[5065]  = 255;
  ram[5066]  = 255;
  ram[5067]  = 255;
  ram[5068]  = 231;
  ram[5069]  = 0;
  ram[5070]  = 190;
  ram[5071]  = 255;
  ram[5072]  = 66;
  ram[5073]  = 42;
  ram[5074]  = 255;
  ram[5075]  = 255;
  ram[5076]  = 255;
  ram[5077]  = 228;
  ram[5078]  = 0;
  ram[5079]  = 208;
  ram[5080]  = 255;
  ram[5081]  = 254;
  ram[5082]  = 255;
  ram[5083]  = 255;
  ram[5084]  = 255;
  ram[5085]  = 143;
  ram[5086]  = 0;
  ram[5087]  = 236;
  ram[5088]  = 255;
  ram[5089]  = 254;
  ram[5090]  = 255;
  ram[5091]  = 120;
  ram[5092]  = 0;
  ram[5093]  = 255;
  ram[5094]  = 249;
  ram[5095]  = 0;
  ram[5096]  = 172;
  ram[5097]  = 255;
  ram[5098]  = 255;
  ram[5099]  = 255;
  ram[5100]  = 58;
  ram[5101]  = 40;
  ram[5102]  = 255;
  ram[5103]  = 255;
  ram[5104]  = 179;
  ram[5105]  = 0;
  ram[5106]  = 245;
  ram[5107]  = 255;
  ram[5108]  = 254;
  ram[5109]  = 255;
  ram[5110]  = 49;
  ram[5111]  = 48;
  ram[5112]  = 255;
  ram[5113]  = 255;
  ram[5114]  = 255;
  ram[5115]  = 0;
  ram[5116]  = 136;
  ram[5117]  = 255;
  ram[5118]  = 252;
  ram[5119]  = 254;
  ram[5120]  = 255;
  ram[5121]  = 35;
  ram[5122]  = 56;
  ram[5123]  = 255;
  ram[5124]  = 227;
  ram[5125]  = 0;
  ram[5126]  = 178;
  ram[5127]  = 255;
  ram[5128]  = 252;
  ram[5129]  = 255;
  ram[5130]  = 28;
  ram[5131]  = 75;
  ram[5132]  = 255;
  ram[5133]  = 254;
  ram[5134]  = 255;
  ram[5135]  = 255;
  ram[5136]  = 254;
  ram[5137]  = 255;
  ram[5138]  = 242;
  ram[5139]  = 0;
  ram[5140]  = 168;
  ram[5141]  = 255;
  ram[5142]  = 255;
  ram[5143]  = 172;
  ram[5144]  = 0;
  ram[5145]  = 237;
  ram[5146]  = 255;
  ram[5147]  = 254;
  ram[5148]  = 255;
  ram[5149]  = 237;
  ram[5150]  = 0;
  ram[5151]  = 165;
  ram[5152]  = 255;
  ram[5153]  = 254;
  ram[5154]  = 255;
  ram[5155]  = 255;
  ram[5156]  = 255;
  ram[5157]  = 147;
  ram[5158]  = 0;
  ram[5159]  = 188;
  ram[5160]  = 255;
  ram[5161]  = 255;
  ram[5162]  = 253;
  ram[5163]  = 252;
  ram[5164]  = 255;
  ram[5165]  = 49;
  ram[5166]  = 49;
  ram[5167]  = 255;
  ram[5168]  = 252;
  ram[5169]  = 251;
  ram[5170]  = 255;
  ram[5171]  = 255;
  ram[5172]  = 255;
  ram[5173]  = 253;
  ram[5174]  = 185;
  ram[5175]  = 0;
  ram[5176]  = 201;
  ram[5177]  = 255;
  ram[5178]  = 161;
  ram[5179]  = 0;
  ram[5180]  = 212;
  ram[5181]  = 255;
  ram[5182]  = 254;
  ram[5183]  = 255;
  ram[5184]  = 207;
  ram[5185]  = 0;
  ram[5186]  = 209;
  ram[5187]  = 255;
  ram[5188]  = 255;
  ram[5189]  = 255;
  ram[5190]  = 255;
  ram[5191]  = 255;
  ram[5192]  = 255;
  ram[5193]  = 255;
  ram[5194]  = 255;
  ram[5195]  = 255;
  ram[5196]  = 235;
  ram[5197]  = 212;
  ram[5198]  = 243;
  ram[5199]  = 255;
  ram[5200]  = 253;
  ram[5201]  = 235;
  ram[5202]  = 209;
  ram[5203]  = 242;
  ram[5204]  = 255;
  ram[5205]  = 254;
  ram[5206]  = 252;
  ram[5207]  = 255;
  ram[5208]  = 255;
  ram[5209]  = 255;
  ram[5210]  = 255;
  ram[5211]  = 255;
  ram[5212]  = 255;
  ram[5213]  = 255;
  ram[5214]  = 255;
  ram[5215]  = 255;
  ram[5216]  = 172;
  ram[5217]  = 0;
  ram[5218]  = 22;
  ram[5219]  = 16;
  ram[5220]  = 29;
  ram[5221]  = 132;
  ram[5222]  = 255;
  ram[5223]  = 252;
  ram[5224]  = 255;
  ram[5225]  = 154;
  ram[5226]  = 0;
  ram[5227]  = 249;
  ram[5228]  = 255;
  ram[5229]  = 255;
  ram[5230]  = 191;
  ram[5231]  = 0;
  ram[5232]  = 23;
  ram[5233]  = 21;
  ram[5234]  = 21;
  ram[5235]  = 23;
  ram[5236]  = 0;
  ram[5237]  = 24;
  ram[5238]  = 255;
  ram[5239]  = 198;
  ram[5240]  = 0;
  ram[5241]  = 0;
  ram[5242]  = 134;
  ram[5243]  = 255;
  ram[5244]  = 255;
  ram[5245]  = 255;
  ram[5246]  = 176;
  ram[5247]  = 0;
  ram[5248]  = 0;
  ram[5249]  = 144;
  ram[5250]  = 255;
  ram[5251]  = 255;
  ram[5252]  = 254;
  ram[5253]  = 253;
  ram[5254]  = 255;
  ram[5255]  = 255;
  ram[5256]  = 255;
  ram[5257]  = 255;
  ram[5258]  = 86;
  ram[5259]  = 8;
  ram[5260]  = 255;
  ram[5261]  = 255;
  ram[5262]  = 255;
  ram[5263]  = 118;
  ram[5264]  = 2;
  ram[5265]  = 255;
  ram[5266]  = 255;
  ram[5267]  = 255;
  ram[5268]  = 234;
  ram[5269]  = 0;
  ram[5270]  = 191;
  ram[5271]  = 255;
  ram[5272]  = 36;
  ram[5273]  = 2;
  ram[5274]  = 24;
  ram[5275]  = 20;
  ram[5276]  = 20;
  ram[5277]  = 20;
  ram[5278]  = 0;
  ram[5279]  = 181;
  ram[5280]  = 255;
  ram[5281]  = 254;
  ram[5282]  = 255;
  ram[5283]  = 255;
  ram[5284]  = 255;
  ram[5285]  = 141;
  ram[5286]  = 0;
  ram[5287]  = 255;
  ram[5288]  = 255;
  ram[5289]  = 254;
  ram[5290]  = 255;
  ram[5291]  = 150;
  ram[5292]  = 0;
  ram[5293]  = 255;
  ram[5294]  = 249;
  ram[5295]  = 0;
  ram[5296]  = 173;
  ram[5297]  = 255;
  ram[5298]  = 255;
  ram[5299]  = 255;
  ram[5300]  = 58;
  ram[5301]  = 41;
  ram[5302]  = 255;
  ram[5303]  = 255;
  ram[5304]  = 180;
  ram[5305]  = 0;
  ram[5306]  = 245;
  ram[5307]  = 255;
  ram[5308]  = 255;
  ram[5309]  = 255;
  ram[5310]  = 50;
  ram[5311]  = 49;
  ram[5312]  = 255;
  ram[5313]  = 255;
  ram[5314]  = 235;
  ram[5315]  = 0;
  ram[5316]  = 184;
  ram[5317]  = 255;
  ram[5318]  = 253;
  ram[5319]  = 253;
  ram[5320]  = 255;
  ram[5321]  = 79;
  ram[5322]  = 17;
  ram[5323]  = 255;
  ram[5324]  = 226;
  ram[5325]  = 0;
  ram[5326]  = 191;
  ram[5327]  = 255;
  ram[5328]  = 255;
  ram[5329]  = 255;
  ram[5330]  = 46;
  ram[5331]  = 72;
  ram[5332]  = 255;
  ram[5333]  = 255;
  ram[5334]  = 255;
  ram[5335]  = 255;
  ram[5336]  = 255;
  ram[5337]  = 255;
  ram[5338]  = 243;
  ram[5339]  = 0;
  ram[5340]  = 168;
  ram[5341]  = 255;
  ram[5342]  = 255;
  ram[5343]  = 121;
  ram[5344]  = 0;
  ram[5345]  = 255;
  ram[5346]  = 255;
  ram[5347]  = 255;
  ram[5348]  = 255;
  ram[5349]  = 255;
  ram[5350]  = 0;
  ram[5351]  = 126;
  ram[5352]  = 255;
  ram[5353]  = 253;
  ram[5354]  = 255;
  ram[5355]  = 255;
  ram[5356]  = 254;
  ram[5357]  = 245;
  ram[5358]  = 0;
  ram[5359]  = 0;
  ram[5360]  = 87;
  ram[5361]  = 249;
  ram[5362]  = 255;
  ram[5363]  = 252;
  ram[5364]  = 255;
  ram[5365]  = 49;
  ram[5366]  = 49;
  ram[5367]  = 255;
  ram[5368]  = 254;
  ram[5369]  = 255;
  ram[5370]  = 255;
  ram[5371]  = 111;
  ram[5372]  = 24;
  ram[5373]  = 0;
  ram[5374]  = 0;
  ram[5375]  = 0;
  ram[5376]  = 203;
  ram[5377]  = 255;
  ram[5378]  = 159;
  ram[5379]  = 0;
  ram[5380]  = 244;
  ram[5381]  = 255;
  ram[5382]  = 255;
  ram[5383]  = 255;
  ram[5384]  = 208;
  ram[5385]  = 0;
  ram[5386]  = 209;
  ram[5387]  = 255;
  ram[5388]  = 255;
  ram[5389]  = 255;
  ram[5390]  = 255;
  ram[5391]  = 255;
  ram[5392]  = 255;
  ram[5393]  = 255;
  ram[5394]  = 255;
  ram[5395]  = 255;
  ram[5396]  = 235;
  ram[5397]  = 212;
  ram[5398]  = 243;
  ram[5399]  = 255;
  ram[5400]  = 253;
  ram[5401]  = 235;
  ram[5402]  = 209;
  ram[5403]  = 242;
  ram[5404]  = 255;
  ram[5405]  = 254;
  ram[5406]  = 252;
  ram[5407]  = 255;
  ram[5408]  = 255;
  ram[5409]  = 255;
  ram[5410]  = 255;
  ram[5411]  = 255;
  ram[5412]  = 255;
  ram[5413]  = 255;
  ram[5414]  = 255;
  ram[5415]  = 255;
  ram[5416]  = 170;
  ram[5417]  = 0;
  ram[5418]  = 238;
  ram[5419]  = 255;
  ram[5420]  = 255;
  ram[5421]  = 255;
  ram[5422]  = 252;
  ram[5423]  = 251;
  ram[5424]  = 255;
  ram[5425]  = 154;
  ram[5426]  = 0;
  ram[5427]  = 247;
  ram[5428]  = 255;
  ram[5429]  = 255;
  ram[5430]  = 187;
  ram[5431]  = 0;
  ram[5432]  = 81;
  ram[5433]  = 89;
  ram[5434]  = 85;
  ram[5435]  = 87;
  ram[5436]  = 85;
  ram[5437]  = 111;
  ram[5438]  = 255;
  ram[5439]  = 255;
  ram[5440]  = 208;
  ram[5441]  = 44;
  ram[5442]  = 0;
  ram[5443]  = 24;
  ram[5444]  = 240;
  ram[5445]  = 255;
  ram[5446]  = 255;
  ram[5447]  = 190;
  ram[5448]  = 28;
  ram[5449]  = 0;
  ram[5450]  = 36;
  ram[5451]  = 255;
  ram[5452]  = 255;
  ram[5453]  = 253;
  ram[5454]  = 255;
  ram[5455]  = 255;
  ram[5456]  = 255;
  ram[5457]  = 255;
  ram[5458]  = 86;
  ram[5459]  = 8;
  ram[5460]  = 255;
  ram[5461]  = 255;
  ram[5462]  = 255;
  ram[5463]  = 118;
  ram[5464]  = 0;
  ram[5465]  = 255;
  ram[5466]  = 255;
  ram[5467]  = 255;
  ram[5468]  = 235;
  ram[5469]  = 0;
  ram[5470]  = 191;
  ram[5471]  = 255;
  ram[5472]  = 30;
  ram[5473]  = 22;
  ram[5474]  = 94;
  ram[5475]  = 86;
  ram[5476]  = 87;
  ram[5477]  = 86;
  ram[5478]  = 81;
  ram[5479]  = 209;
  ram[5480]  = 255;
  ram[5481]  = 254;
  ram[5482]  = 255;
  ram[5483]  = 255;
  ram[5484]  = 255;
  ram[5485]  = 141;
  ram[5486]  = 0;
  ram[5487]  = 255;
  ram[5488]  = 253;
  ram[5489]  = 254;
  ram[5490]  = 255;
  ram[5491]  = 147;
  ram[5492]  = 0;
  ram[5493]  = 255;
  ram[5494]  = 248;
  ram[5495]  = 0;
  ram[5496]  = 174;
  ram[5497]  = 255;
  ram[5498]  = 255;
  ram[5499]  = 255;
  ram[5500]  = 60;
  ram[5501]  = 40;
  ram[5502]  = 255;
  ram[5503]  = 255;
  ram[5504]  = 179;
  ram[5505]  = 0;
  ram[5506]  = 246;
  ram[5507]  = 255;
  ram[5508]  = 255;
  ram[5509]  = 255;
  ram[5510]  = 50;
  ram[5511]  = 49;
  ram[5512]  = 255;
  ram[5513]  = 255;
  ram[5514]  = 230;
  ram[5515]  = 0;
  ram[5516]  = 190;
  ram[5517]  = 255;
  ram[5518]  = 254;
  ram[5519]  = 254;
  ram[5520]  = 255;
  ram[5521]  = 83;
  ram[5522]  = 18;
  ram[5523]  = 255;
  ram[5524]  = 227;
  ram[5525]  = 0;
  ram[5526]  = 191;
  ram[5527]  = 255;
  ram[5528]  = 254;
  ram[5529]  = 255;
  ram[5530]  = 47;
  ram[5531]  = 72;
  ram[5532]  = 255;
  ram[5533]  = 255;
  ram[5534]  = 255;
  ram[5535]  = 255;
  ram[5536]  = 255;
  ram[5537]  = 255;
  ram[5538]  = 242;
  ram[5539]  = 0;
  ram[5540]  = 168;
  ram[5541]  = 255;
  ram[5542]  = 255;
  ram[5543]  = 119;
  ram[5544]  = 0;
  ram[5545]  = 255;
  ram[5546]  = 255;
  ram[5547]  = 255;
  ram[5548]  = 255;
  ram[5549]  = 255;
  ram[5550]  = 0;
  ram[5551]  = 126;
  ram[5552]  = 255;
  ram[5553]  = 254;
  ram[5554]  = 255;
  ram[5555]  = 255;
  ram[5556]  = 253;
  ram[5557]  = 255;
  ram[5558]  = 240;
  ram[5559]  = 70;
  ram[5560]  = 0;
  ram[5561]  = 0;
  ram[5562]  = 207;
  ram[5563]  = 255;
  ram[5564]  = 255;
  ram[5565]  = 49;
  ram[5566]  = 49;
  ram[5567]  = 255;
  ram[5568]  = 253;
  ram[5569]  = 255;
  ram[5570]  = 58;
  ram[5571]  = 0;
  ram[5572]  = 100;
  ram[5573]  = 170;
  ram[5574]  = 205;
  ram[5575]  = 0;
  ram[5576]  = 202;
  ram[5577]  = 255;
  ram[5578]  = 159;
  ram[5579]  = 0;
  ram[5580]  = 243;
  ram[5581]  = 255;
  ram[5582]  = 255;
  ram[5583]  = 255;
  ram[5584]  = 208;
  ram[5585]  = 0;
  ram[5586]  = 209;
  ram[5587]  = 255;
  ram[5588]  = 255;
  ram[5589]  = 255;
  ram[5590]  = 255;
  ram[5591]  = 255;
  ram[5592]  = 255;
  ram[5593]  = 255;
  ram[5594]  = 255;
  ram[5595]  = 255;
  ram[5596]  = 236;
  ram[5597]  = 211;
  ram[5598]  = 243;
  ram[5599]  = 255;
  ram[5600]  = 253;
  ram[5601]  = 235;
  ram[5602]  = 209;
  ram[5603]  = 242;
  ram[5604]  = 255;
  ram[5605]  = 254;
  ram[5606]  = 252;
  ram[5607]  = 255;
  ram[5608]  = 255;
  ram[5609]  = 255;
  ram[5610]  = 255;
  ram[5611]  = 255;
  ram[5612]  = 255;
  ram[5613]  = 255;
  ram[5614]  = 255;
  ram[5615]  = 255;
  ram[5616]  = 170;
  ram[5617]  = 0;
  ram[5618]  = 230;
  ram[5619]  = 255;
  ram[5620]  = 255;
  ram[5621]  = 253;
  ram[5622]  = 253;
  ram[5623]  = 254;
  ram[5624]  = 255;
  ram[5625]  = 153;
  ram[5626]  = 0;
  ram[5627]  = 248;
  ram[5628]  = 255;
  ram[5629]  = 255;
  ram[5630]  = 208;
  ram[5631]  = 0;
  ram[5632]  = 218;
  ram[5633]  = 255;
  ram[5634]  = 255;
  ram[5635]  = 255;
  ram[5636]  = 255;
  ram[5637]  = 255;
  ram[5638]  = 254;
  ram[5639]  = 252;
  ram[5640]  = 255;
  ram[5641]  = 255;
  ram[5642]  = 147;
  ram[5643]  = 0;
  ram[5644]  = 118;
  ram[5645]  = 255;
  ram[5646]  = 253;
  ram[5647]  = 255;
  ram[5648]  = 253;
  ram[5649]  = 126;
  ram[5650]  = 0;
  ram[5651]  = 150;
  ram[5652]  = 255;
  ram[5653]  = 253;
  ram[5654]  = 253;
  ram[5655]  = 253;
  ram[5656]  = 253;
  ram[5657]  = 255;
  ram[5658]  = 87;
  ram[5659]  = 9;
  ram[5660]  = 255;
  ram[5661]  = 252;
  ram[5662]  = 255;
  ram[5663]  = 120;
  ram[5664]  = 0;
  ram[5665]  = 255;
  ram[5666]  = 255;
  ram[5667]  = 255;
  ram[5668]  = 234;
  ram[5669]  = 0;
  ram[5670]  = 191;
  ram[5671]  = 255;
  ram[5672]  = 38;
  ram[5673]  = 59;
  ram[5674]  = 255;
  ram[5675]  = 255;
  ram[5676]  = 255;
  ram[5677]  = 255;
  ram[5678]  = 255;
  ram[5679]  = 255;
  ram[5680]  = 255;
  ram[5681]  = 255;
  ram[5682]  = 255;
  ram[5683]  = 255;
  ram[5684]  = 255;
  ram[5685]  = 141;
  ram[5686]  = 0;
  ram[5687]  = 255;
  ram[5688]  = 255;
  ram[5689]  = 252;
  ram[5690]  = 255;
  ram[5691]  = 118;
  ram[5692]  = 0;
  ram[5693]  = 255;
  ram[5694]  = 248;
  ram[5695]  = 0;
  ram[5696]  = 169;
  ram[5697]  = 255;
  ram[5698]  = 254;
  ram[5699]  = 255;
  ram[5700]  = 52;
  ram[5701]  = 41;
  ram[5702]  = 255;
  ram[5703]  = 255;
  ram[5704]  = 180;
  ram[5705]  = 0;
  ram[5706]  = 246;
  ram[5707]  = 255;
  ram[5708]  = 254;
  ram[5709]  = 255;
  ram[5710]  = 50;
  ram[5711]  = 48;
  ram[5712]  = 255;
  ram[5713]  = 255;
  ram[5714]  = 245;
  ram[5715]  = 0;
  ram[5716]  = 163;
  ram[5717]  = 255;
  ram[5718]  = 252;
  ram[5719]  = 252;
  ram[5720]  = 255;
  ram[5721]  = 61;
  ram[5722]  = 43;
  ram[5723]  = 255;
  ram[5724]  = 225;
  ram[5725]  = 0;
  ram[5726]  = 191;
  ram[5727]  = 255;
  ram[5728]  = 254;
  ram[5729]  = 255;
  ram[5730]  = 46;
  ram[5731]  = 72;
  ram[5732]  = 255;
  ram[5733]  = 255;
  ram[5734]  = 255;
  ram[5735]  = 255;
  ram[5736]  = 255;
  ram[5737]  = 255;
  ram[5738]  = 243;
  ram[5739]  = 0;
  ram[5740]  = 168;
  ram[5741]  = 255;
  ram[5742]  = 255;
  ram[5743]  = 143;
  ram[5744]  = 0;
  ram[5745]  = 255;
  ram[5746]  = 255;
  ram[5747]  = 253;
  ram[5748]  = 255;
  ram[5749]  = 252;
  ram[5750]  = 0;
  ram[5751]  = 154;
  ram[5752]  = 255;
  ram[5753]  = 253;
  ram[5754]  = 255;
  ram[5755]  = 255;
  ram[5756]  = 251;
  ram[5757]  = 251;
  ram[5758]  = 255;
  ram[5759]  = 255;
  ram[5760]  = 187;
  ram[5761]  = 0;
  ram[5762]  = 51;
  ram[5763]  = 255;
  ram[5764]  = 255;
  ram[5765]  = 49;
  ram[5766]  = 49;
  ram[5767]  = 255;
  ram[5768]  = 255;
  ram[5769]  = 237;
  ram[5770]  = 0;
  ram[5771]  = 152;
  ram[5772]  = 255;
  ram[5773]  = 255;
  ram[5774]  = 229;
  ram[5775]  = 0;
  ram[5776]  = 202;
  ram[5777]  = 255;
  ram[5778]  = 158;
  ram[5779]  = 0;
  ram[5780]  = 244;
  ram[5781]  = 255;
  ram[5782]  = 255;
  ram[5783]  = 255;
  ram[5784]  = 208;
  ram[5785]  = 0;
  ram[5786]  = 210;
  ram[5787]  = 255;
  ram[5788]  = 255;
  ram[5789]  = 255;
  ram[5790]  = 255;
  ram[5791]  = 255;
  ram[5792]  = 255;
  ram[5793]  = 255;
  ram[5794]  = 255;
  ram[5795]  = 255;
  ram[5796]  = 236;
  ram[5797]  = 211;
  ram[5798]  = 243;
  ram[5799]  = 255;
  ram[5800]  = 253;
  ram[5801]  = 235;
  ram[5802]  = 209;
  ram[5803]  = 242;
  ram[5804]  = 255;
  ram[5805]  = 254;
  ram[5806]  = 252;
  ram[5807]  = 255;
  ram[5808]  = 255;
  ram[5809]  = 255;
  ram[5810]  = 255;
  ram[5811]  = 255;
  ram[5812]  = 255;
  ram[5813]  = 255;
  ram[5814]  = 255;
  ram[5815]  = 255;
  ram[5816]  = 170;
  ram[5817]  = 0;
  ram[5818]  = 230;
  ram[5819]  = 255;
  ram[5820]  = 255;
  ram[5821]  = 255;
  ram[5822]  = 255;
  ram[5823]  = 255;
  ram[5824]  = 255;
  ram[5825]  = 153;
  ram[5826]  = 0;
  ram[5827]  = 250;
  ram[5828]  = 255;
  ram[5829]  = 255;
  ram[5830]  = 243;
  ram[5831]  = 0;
  ram[5832]  = 135;
  ram[5833]  = 255;
  ram[5834]  = 253;
  ram[5835]  = 255;
  ram[5836]  = 255;
  ram[5837]  = 255;
  ram[5838]  = 254;
  ram[5839]  = 255;
  ram[5840]  = 255;
  ram[5841]  = 255;
  ram[5842]  = 255;
  ram[5843]  = 36;
  ram[5844]  = 65;
  ram[5845]  = 255;
  ram[5846]  = 255;
  ram[5847]  = 255;
  ram[5848]  = 255;
  ram[5849]  = 255;
  ram[5850]  = 13;
  ram[5851]  = 84;
  ram[5852]  = 255;
  ram[5853]  = 252;
  ram[5854]  = 252;
  ram[5855]  = 253;
  ram[5856]  = 253;
  ram[5857]  = 255;
  ram[5858]  = 86;
  ram[5859]  = 13;
  ram[5860]  = 255;
  ram[5861]  = 255;
  ram[5862]  = 255;
  ram[5863]  = 118;
  ram[5864]  = 0;
  ram[5865]  = 255;
  ram[5866]  = 255;
  ram[5867]  = 255;
  ram[5868]  = 234;
  ram[5869]  = 0;
  ram[5870]  = 191;
  ram[5871]  = 255;
  ram[5872]  = 92;
  ram[5873]  = 0;
  ram[5874]  = 255;
  ram[5875]  = 255;
  ram[5876]  = 251;
  ram[5877]  = 255;
  ram[5878]  = 255;
  ram[5879]  = 255;
  ram[5880]  = 255;
  ram[5881]  = 255;
  ram[5882]  = 255;
  ram[5883]  = 255;
  ram[5884]  = 255;
  ram[5885]  = 144;
  ram[5886]  = 0;
  ram[5887]  = 217;
  ram[5888]  = 255;
  ram[5889]  = 254;
  ram[5890]  = 255;
  ram[5891]  = 32;
  ram[5892]  = 38;
  ram[5893]  = 255;
  ram[5894]  = 248;
  ram[5895]  = 0;
  ram[5896]  = 128;
  ram[5897]  = 255;
  ram[5898]  = 251;
  ram[5899]  = 255;
  ram[5900]  = 12;
  ram[5901]  = 45;
  ram[5902]  = 255;
  ram[5903]  = 255;
  ram[5904]  = 179;
  ram[5905]  = 0;
  ram[5906]  = 253;
  ram[5907]  = 255;
  ram[5908]  = 252;
  ram[5909]  = 255;
  ram[5910]  = 44;
  ram[5911]  = 52;
  ram[5912]  = 255;
  ram[5913]  = 253;
  ram[5914]  = 255;
  ram[5915]  = 0;
  ram[5916]  = 72;
  ram[5917]  = 255;
  ram[5918]  = 255;
  ram[5919]  = 255;
  ram[5920]  = 255;
  ram[5921]  = 0;
  ram[5922]  = 115;
  ram[5923]  = 255;
  ram[5924]  = 225;
  ram[5925]  = 0;
  ram[5926]  = 191;
  ram[5927]  = 255;
  ram[5928]  = 255;
  ram[5929]  = 255;
  ram[5930]  = 47;
  ram[5931]  = 72;
  ram[5932]  = 255;
  ram[5933]  = 255;
  ram[5934]  = 255;
  ram[5935]  = 255;
  ram[5936]  = 255;
  ram[5937]  = 255;
  ram[5938]  = 241;
  ram[5939]  = 0;
  ram[5940]  = 175;
  ram[5941]  = 255;
  ram[5942]  = 255;
  ram[5943]  = 202;
  ram[5944]  = 0;
  ram[5945]  = 182;
  ram[5946]  = 255;
  ram[5947]  = 255;
  ram[5948]  = 255;
  ram[5949]  = 197;
  ram[5950]  = 0;
  ram[5951]  = 214;
  ram[5952]  = 255;
  ram[5953]  = 253;
  ram[5954]  = 255;
  ram[5955]  = 255;
  ram[5956]  = 254;
  ram[5957]  = 255;
  ram[5958]  = 255;
  ram[5959]  = 255;
  ram[5960]  = 255;
  ram[5961]  = 107;
  ram[5962]  = 0;
  ram[5963]  = 255;
  ram[5964]  = 255;
  ram[5965]  = 45;
  ram[5966]  = 54;
  ram[5967]  = 255;
  ram[5968]  = 255;
  ram[5969]  = 213;
  ram[5970]  = 0;
  ram[5971]  = 224;
  ram[5972]  = 255;
  ram[5973]  = 255;
  ram[5974]  = 179;
  ram[5975]  = 0;
  ram[5976]  = 201;
  ram[5977]  = 255;
  ram[5978]  = 158;
  ram[5979]  = 0;
  ram[5980]  = 244;
  ram[5981]  = 255;
  ram[5982]  = 255;
  ram[5983]  = 255;
  ram[5984]  = 204;
  ram[5985]  = 0;
  ram[5986]  = 215;
  ram[5987]  = 255;
  ram[5988]  = 252;
  ram[5989]  = 255;
  ram[5990]  = 255;
  ram[5991]  = 255;
  ram[5992]  = 255;
  ram[5993]  = 255;
  ram[5994]  = 255;
  ram[5995]  = 255;
  ram[5996]  = 236;
  ram[5997]  = 211;
  ram[5998]  = 243;
  ram[5999]  = 255;
  ram[6000]  = 253;
  ram[6001]  = 235;
  ram[6002]  = 209;
  ram[6003]  = 242;
  ram[6004]  = 255;
  ram[6005]  = 254;
  ram[6006]  = 252;
  ram[6007]  = 255;
  ram[6008]  = 255;
  ram[6009]  = 255;
  ram[6010]  = 255;
  ram[6011]  = 255;
  ram[6012]  = 255;
  ram[6013]  = 255;
  ram[6014]  = 255;
  ram[6015]  = 255;
  ram[6016]  = 170;
  ram[6017]  = 0;
  ram[6018]  = 230;
  ram[6019]  = 255;
  ram[6020]  = 255;
  ram[6021]  = 255;
  ram[6022]  = 255;
  ram[6023]  = 255;
  ram[6024]  = 255;
  ram[6025]  = 153;
  ram[6026]  = 0;
  ram[6027]  = 250;
  ram[6028]  = 255;
  ram[6029]  = 254;
  ram[6030]  = 255;
  ram[6031]  = 64;
  ram[6032]  = 0;
  ram[6033]  = 204;
  ram[6034]  = 255;
  ram[6035]  = 255;
  ram[6036]  = 127;
  ram[6037]  = 208;
  ram[6038]  = 255;
  ram[6039]  = 135;
  ram[6040]  = 234;
  ram[6041]  = 255;
  ram[6042]  = 252;
  ram[6043]  = 0;
  ram[6044]  = 97;
  ram[6045]  = 255;
  ram[6046]  = 120;
  ram[6047]  = 244;
  ram[6048]  = 255;
  ram[6049]  = 233;
  ram[6050]  = 0;
  ram[6051]  = 125;
  ram[6052]  = 255;
  ram[6053]  = 255;
  ram[6054]  = 254;
  ram[6055]  = 254;
  ram[6056]  = 253;
  ram[6057]  = 255;
  ram[6058]  = 112;
  ram[6059]  = 0;
  ram[6060]  = 243;
  ram[6061]  = 245;
  ram[6062]  = 255;
  ram[6063]  = 120;
  ram[6064]  = 0;
  ram[6065]  = 255;
  ram[6066]  = 255;
  ram[6067]  = 255;
  ram[6068]  = 234;
  ram[6069]  = 0;
  ram[6070]  = 191;
  ram[6071]  = 255;
  ram[6072]  = 212;
  ram[6073]  = 0;
  ram[6074]  = 92;
  ram[6075]  = 255;
  ram[6076]  = 255;
  ram[6077]  = 215;
  ram[6078]  = 114;
  ram[6079]  = 255;
  ram[6080]  = 255;
  ram[6081]  = 255;
  ram[6082]  = 255;
  ram[6083]  = 255;
  ram[6084]  = 255;
  ram[6085]  = 145;
  ram[6086]  = 0;
  ram[6087]  = 39;
  ram[6088]  = 243;
  ram[6089]  = 255;
  ram[6090]  = 134;
  ram[6091]  = 0;
  ram[6092]  = 174;
  ram[6093]  = 255;
  ram[6094]  = 255;
  ram[6095]  = 39;
  ram[6096]  = 2;
  ram[6097]  = 237;
  ram[6098]  = 255;
  ram[6099]  = 117;
  ram[6100]  = 0;
  ram[6101]  = 50;
  ram[6102]  = 255;
  ram[6103]  = 255;
  ram[6104]  = 202;
  ram[6105]  = 0;
  ram[6106]  = 173;
  ram[6107]  = 255;
  ram[6108]  = 249;
  ram[6109]  = 255;
  ram[6110]  = 78;
  ram[6111]  = 8;
  ram[6112]  = 255;
  ram[6113]  = 245;
  ram[6114]  = 255;
  ram[6115]  = 130;
  ram[6116]  = 0;
  ram[6117]  = 156;
  ram[6118]  = 255;
  ram[6119]  = 255;
  ram[6120]  = 90;
  ram[6121]  = 0;
  ram[6122]  = 234;
  ram[6123]  = 255;
  ram[6124]  = 225;
  ram[6125]  = 0;
  ram[6126]  = 191;
  ram[6127]  = 255;
  ram[6128]  = 255;
  ram[6129]  = 255;
  ram[6130]  = 47;
  ram[6131]  = 72;
  ram[6132]  = 255;
  ram[6133]  = 255;
  ram[6134]  = 255;
  ram[6135]  = 255;
  ram[6136]  = 255;
  ram[6137]  = 255;
  ram[6138]  = 255;
  ram[6139]  = 0;
  ram[6140]  = 94;
  ram[6141]  = 255;
  ram[6142]  = 246;
  ram[6143]  = 255;
  ram[6144]  = 21;
  ram[6145]  = 0;
  ram[6146]  = 224;
  ram[6147]  = 255;
  ram[6148]  = 239;
  ram[6149]  = 3;
  ram[6150]  = 44;
  ram[6151]  = 255;
  ram[6152]  = 254;
  ram[6153]  = 254;
  ram[6154]  = 255;
  ram[6155]  = 255;
  ram[6156]  = 255;
  ram[6157]  = 156;
  ram[6158]  = 209;
  ram[6159]  = 255;
  ram[6160]  = 255;
  ram[6161]  = 44;
  ram[6162]  = 30;
  ram[6163]  = 255;
  ram[6164]  = 255;
  ram[6165]  = 79;
  ram[6166]  = 10;
  ram[6167]  = 255;
  ram[6168]  = 250;
  ram[6169]  = 234;
  ram[6170]  = 0;
  ram[6171]  = 114;
  ram[6172]  = 255;
  ram[6173]  = 238;
  ram[6174]  = 7;
  ram[6175]  = 0;
  ram[6176]  = 203;
  ram[6177]  = 255;
  ram[6178]  = 158;
  ram[6179]  = 0;
  ram[6180]  = 244;
  ram[6181]  = 255;
  ram[6182]  = 255;
  ram[6183]  = 255;
  ram[6184]  = 225;
  ram[6185]  = 0;
  ram[6186]  = 148;
  ram[6187]  = 255;
  ram[6188]  = 248;
  ram[6189]  = 255;
  ram[6190]  = 255;
  ram[6191]  = 255;
  ram[6192]  = 255;
  ram[6193]  = 255;
  ram[6194]  = 255;
  ram[6195]  = 255;
  ram[6196]  = 236;
  ram[6197]  = 211;
  ram[6198]  = 243;
  ram[6199]  = 255;
  ram[6200]  = 253;
  ram[6201]  = 235;
  ram[6202]  = 209;
  ram[6203]  = 242;
  ram[6204]  = 255;
  ram[6205]  = 254;
  ram[6206]  = 252;
  ram[6207]  = 255;
  ram[6208]  = 255;
  ram[6209]  = 255;
  ram[6210]  = 255;
  ram[6211]  = 255;
  ram[6212]  = 255;
  ram[6213]  = 255;
  ram[6214]  = 253;
  ram[6215]  = 255;
  ram[6216]  = 164;
  ram[6217]  = 0;
  ram[6218]  = 226;
  ram[6219]  = 255;
  ram[6220]  = 255;
  ram[6221]  = 255;
  ram[6222]  = 255;
  ram[6223]  = 255;
  ram[6224]  = 255;
  ram[6225]  = 144;
  ram[6226]  = 0;
  ram[6227]  = 247;
  ram[6228]  = 255;
  ram[6229]  = 251;
  ram[6230]  = 255;
  ram[6231]  = 222;
  ram[6232]  = 1;
  ram[6233]  = 0;
  ram[6234]  = 32;
  ram[6235]  = 10;
  ram[6236]  = 0;
  ram[6237]  = 220;
  ram[6238]  = 255;
  ram[6239]  = 41;
  ram[6240]  = 0;
  ram[6241]  = 31;
  ram[6242]  = 1;
  ram[6243]  = 0;
  ram[6244]  = 221;
  ram[6245]  = 255;
  ram[6246]  = 7;
  ram[6247]  = 0;
  ram[6248]  = 30;
  ram[6249]  = 0;
  ram[6250]  = 6;
  ram[6251]  = 246;
  ram[6252]  = 255;
  ram[6253]  = 254;
  ram[6254]  = 255;
  ram[6255]  = 255;
  ram[6256]  = 254;
  ram[6257]  = 255;
  ram[6258]  = 201;
  ram[6259]  = 0;
  ram[6260]  = 0;
  ram[6261]  = 50;
  ram[6262]  = 255;
  ram[6263]  = 110;
  ram[6264]  = 0;
  ram[6265]  = 255;
  ram[6266]  = 254;
  ram[6267]  = 255;
  ram[6268]  = 231;
  ram[6269]  = 0;
  ram[6270]  = 183;
  ram[6271]  = 255;
  ram[6272]  = 255;
  ram[6273]  = 98;
  ram[6274]  = 0;
  ram[6275]  = 14;
  ram[6276]  = 26;
  ram[6277]  = 0;
  ram[6278]  = 77;
  ram[6279]  = 255;
  ram[6280]  = 255;
  ram[6281]  = 255;
  ram[6282]  = 255;
  ram[6283]  = 255;
  ram[6284]  = 255;
  ram[6285]  = 135;
  ram[6286]  = 0;
  ram[6287]  = 70;
  ram[6288]  = 0;
  ram[6289]  = 19;
  ram[6290]  = 0;
  ram[6291]  = 63;
  ram[6292]  = 255;
  ram[6293]  = 253;
  ram[6294]  = 255;
  ram[6295]  = 161;
  ram[6296]  = 0;
  ram[6297]  = 0;
  ram[6298]  = 14;
  ram[6299]  = 47;
  ram[6300]  = 51;
  ram[6301]  = 29;
  ram[6302]  = 255;
  ram[6303]  = 255;
  ram[6304]  = 254;
  ram[6305]  = 10;
  ram[6306]  = 0;
  ram[6307]  = 13;
  ram[6308]  = 225;
  ram[6309]  = 255;
  ram[6310]  = 177;
  ram[6311]  = 0;
  ram[6312]  = 2;
  ram[6313]  = 74;
  ram[6314]  = 255;
  ram[6315]  = 255;
  ram[6316]  = 47;
  ram[6317]  = 0;
  ram[6318]  = 22;
  ram[6319]  = 11;
  ram[6320]  = 0;
  ram[6321]  = 140;
  ram[6322]  = 255;
  ram[6323]  = 255;
  ram[6324]  = 221;
  ram[6325]  = 0;
  ram[6326]  = 185;
  ram[6327]  = 255;
  ram[6328]  = 255;
  ram[6329]  = 255;
  ram[6330]  = 33;
  ram[6331]  = 61;
  ram[6332]  = 255;
  ram[6333]  = 252;
  ram[6334]  = 255;
  ram[6335]  = 255;
  ram[6336]  = 255;
  ram[6337]  = 255;
  ram[6338]  = 255;
  ram[6339]  = 72;
  ram[6340]  = 0;
  ram[6341]  = 4;
  ram[6342]  = 159;
  ram[6343]  = 255;
  ram[6344]  = 217;
  ram[6345]  = 0;
  ram[6346]  = 0;
  ram[6347]  = 24;
  ram[6348]  = 0;
  ram[6349]  = 3;
  ram[6350]  = 217;
  ram[6351]  = 255;
  ram[6352]  = 252;
  ram[6353]  = 253;
  ram[6354]  = 255;
  ram[6355]  = 255;
  ram[6356]  = 255;
  ram[6357]  = 111;
  ram[6358]  = 0;
  ram[6359]  = 28;
  ram[6360]  = 17;
  ram[6361]  = 0;
  ram[6362]  = 176;
  ram[6363]  = 255;
  ram[6364]  = 255;
  ram[6365]  = 175;
  ram[6366]  = 0;
  ram[6367]  = 2;
  ram[6368]  = 77;
  ram[6369]  = 255;
  ram[6370]  = 44;
  ram[6371]  = 0;
  ram[6372]  = 26;
  ram[6373]  = 0;
  ram[6374]  = 133;
  ram[6375]  = 0;
  ram[6376]  = 197;
  ram[6377]  = 255;
  ram[6378]  = 151;
  ram[6379]  = 0;
  ram[6380]  = 242;
  ram[6381]  = 255;
  ram[6382]  = 255;
  ram[6383]  = 255;
  ram[6384]  = 255;
  ram[6385]  = 34;
  ram[6386]  = 0;
  ram[6387]  = 1;
  ram[6388]  = 210;
  ram[6389]  = 255;
  ram[6390]  = 255;
  ram[6391]  = 255;
  ram[6392]  = 255;
  ram[6393]  = 255;
  ram[6394]  = 255;
  ram[6395]  = 255;
  ram[6396]  = 235;
  ram[6397]  = 212;
  ram[6398]  = 243;
  ram[6399]  = 255;
  ram[6400]  = 253;
  ram[6401]  = 235;
  ram[6402]  = 209;
  ram[6403]  = 242;
  ram[6404]  = 255;
  ram[6405]  = 254;
  ram[6406]  = 252;
  ram[6407]  = 255;
  ram[6408]  = 255;
  ram[6409]  = 255;
  ram[6410]  = 255;
  ram[6411]  = 255;
  ram[6412]  = 255;
  ram[6413]  = 255;
  ram[6414]  = 253;
  ram[6415]  = 255;
  ram[6416]  = 213;
  ram[6417]  = 129;
  ram[6418]  = 240;
  ram[6419]  = 255;
  ram[6420]  = 255;
  ram[6421]  = 255;
  ram[6422]  = 255;
  ram[6423]  = 255;
  ram[6424]  = 255;
  ram[6425]  = 206;
  ram[6426]  = 134;
  ram[6427]  = 250;
  ram[6428]  = 253;
  ram[6429]  = 255;
  ram[6430]  = 255;
  ram[6431]  = 255;
  ram[6432]  = 216;
  ram[6433]  = 96;
  ram[6434]  = 50;
  ram[6435]  = 91;
  ram[6436]  = 193;
  ram[6437]  = 255;
  ram[6438]  = 255;
  ram[6439]  = 199;
  ram[6440]  = 92;
  ram[6441]  = 52;
  ram[6442]  = 102;
  ram[6443]  = 223;
  ram[6444]  = 255;
  ram[6445]  = 255;
  ram[6446]  = 184;
  ram[6447]  = 82;
  ram[6448]  = 53;
  ram[6449]  = 109;
  ram[6450]  = 232;
  ram[6451]  = 255;
  ram[6452]  = 255;
  ram[6453]  = 255;
  ram[6454]  = 255;
  ram[6455]  = 255;
  ram[6456]  = 254;
  ram[6457]  = 251;
  ram[6458]  = 255;
  ram[6459]  = 152;
  ram[6460]  = 62;
  ram[6461]  = 133;
  ram[6462]  = 255;
  ram[6463]  = 192;
  ram[6464]  = 139;
  ram[6465]  = 255;
  ram[6466]  = 252;
  ram[6467]  = 253;
  ram[6468]  = 240;
  ram[6469]  = 120;
  ram[6470]  = 218;
  ram[6471]  = 255;
  ram[6472]  = 255;
  ram[6473]  = 255;
  ram[6474]  = 145;
  ram[6475]  = 61;
  ram[6476]  = 67;
  ram[6477]  = 140;
  ram[6478]  = 242;
  ram[6479]  = 255;
  ram[6480]  = 255;
  ram[6481]  = 255;
  ram[6482]  = 255;
  ram[6483]  = 255;
  ram[6484]  = 255;
  ram[6485]  = 200;
  ram[6486]  = 141;
  ram[6487]  = 252;
  ram[6488]  = 116;
  ram[6489]  = 51;
  ram[6490]  = 126;
  ram[6491]  = 250;
  ram[6492]  = 255;
  ram[6493]  = 254;
  ram[6494]  = 250;
  ram[6495]  = 255;
  ram[6496]  = 155;
  ram[6497]  = 56;
  ram[6498]  = 89;
  ram[6499]  = 236;
  ram[6500]  = 175;
  ram[6501]  = 155;
  ram[6502]  = 255;
  ram[6503]  = 251;
  ram[6504]  = 255;
  ram[6505]  = 202;
  ram[6506]  = 70;
  ram[6507]  = 91;
  ram[6508]  = 244;
  ram[6509]  = 254;
  ram[6510]  = 255;
  ram[6511]  = 132;
  ram[6512]  = 60;
  ram[6513]  = 152;
  ram[6514]  = 255;
  ram[6515]  = 255;
  ram[6516]  = 247;
  ram[6517]  = 137;
  ram[6518]  = 61;
  ram[6519]  = 76;
  ram[6520]  = 182;
  ram[6521]  = 255;
  ram[6522]  = 255;
  ram[6523]  = 255;
  ram[6524]  = 237;
  ram[6525]  = 124;
  ram[6526]  = 226;
  ram[6527]  = 255;
  ram[6528]  = 254;
  ram[6529]  = 255;
  ram[6530]  = 160;
  ram[6531]  = 172;
  ram[6532]  = 255;
  ram[6533]  = 252;
  ram[6534]  = 255;
  ram[6535]  = 255;
  ram[6536]  = 255;
  ram[6537]  = 255;
  ram[6538]  = 255;
  ram[6539]  = 239;
  ram[6540]  = 88;
  ram[6541]  = 69;
  ram[6542]  = 209;
  ram[6543]  = 255;
  ram[6544]  = 255;
  ram[6545]  = 216;
  ram[6546]  = 100;
  ram[6547]  = 51;
  ram[6548]  = 102;
  ram[6549]  = 227;
  ram[6550]  = 255;
  ram[6551]  = 255;
  ram[6552]  = 255;
  ram[6553]  = 255;
  ram[6554]  = 255;
  ram[6555]  = 255;
  ram[6556]  = 255;
  ram[6557]  = 224;
  ram[6558]  = 109;
  ram[6559]  = 52;
  ram[6560]  = 83;
  ram[6561]  = 196;
  ram[6562]  = 255;
  ram[6563]  = 253;
  ram[6564]  = 252;
  ram[6565]  = 255;
  ram[6566]  = 131;
  ram[6567]  = 62;
  ram[6568]  = 154;
  ram[6569]  = 255;
  ram[6570]  = 239;
  ram[6571]  = 100;
  ram[6572]  = 51;
  ram[6573]  = 154;
  ram[6574]  = 255;
  ram[6575]  = 124;
  ram[6576]  = 228;
  ram[6577]  = 255;
  ram[6578]  = 211;
  ram[6579]  = 130;
  ram[6580]  = 247;
  ram[6581]  = 255;
  ram[6582]  = 255;
  ram[6583]  = 253;
  ram[6584]  = 255;
  ram[6585]  = 215;
  ram[6586]  = 79;
  ram[6587]  = 76;
  ram[6588]  = 239;
  ram[6589]  = 255;
  ram[6590]  = 255;
  ram[6591]  = 255;
  ram[6592]  = 255;
  ram[6593]  = 255;
  ram[6594]  = 255;
  ram[6595]  = 255;
  ram[6596]  = 236;
  ram[6597]  = 212;
  ram[6598]  = 243;
  ram[6599]  = 255;
  ram[6600]  = 253;
  ram[6601]  = 235;
  ram[6602]  = 209;
  ram[6603]  = 242;
  ram[6604]  = 255;
  ram[6605]  = 254;
  ram[6606]  = 252;
  ram[6607]  = 255;
  ram[6608]  = 255;
  ram[6609]  = 255;
  ram[6610]  = 255;
  ram[6611]  = 255;
  ram[6612]  = 255;
  ram[6613]  = 255;
  ram[6614]  = 254;
  ram[6615]  = 251;
  ram[6616]  = 253;
  ram[6617]  = 255;
  ram[6618]  = 255;
  ram[6619]  = 253;
  ram[6620]  = 255;
  ram[6621]  = 255;
  ram[6622]  = 255;
  ram[6623]  = 255;
  ram[6624]  = 251;
  ram[6625]  = 255;
  ram[6626]  = 255;
  ram[6627]  = 254;
  ram[6628]  = 253;
  ram[6629]  = 253;
  ram[6630]  = 255;
  ram[6631]  = 255;
  ram[6632]  = 255;
  ram[6633]  = 255;
  ram[6634]  = 255;
  ram[6635]  = 255;
  ram[6636]  = 255;
  ram[6637]  = 252;
  ram[6638]  = 252;
  ram[6639]  = 255;
  ram[6640]  = 255;
  ram[6641]  = 255;
  ram[6642]  = 255;
  ram[6643]  = 255;
  ram[6644]  = 250;
  ram[6645]  = 253;
  ram[6646]  = 255;
  ram[6647]  = 255;
  ram[6648]  = 255;
  ram[6649]  = 255;
  ram[6650]  = 255;
  ram[6651]  = 251;
  ram[6652]  = 255;
  ram[6653]  = 255;
  ram[6654]  = 255;
  ram[6655]  = 255;
  ram[6656]  = 254;
  ram[6657]  = 252;
  ram[6658]  = 252;
  ram[6659]  = 255;
  ram[6660]  = 255;
  ram[6661]  = 255;
  ram[6662]  = 254;
  ram[6663]  = 255;
  ram[6664]  = 255;
  ram[6665]  = 253;
  ram[6666]  = 252;
  ram[6667]  = 253;
  ram[6668]  = 251;
  ram[6669]  = 255;
  ram[6670]  = 255;
  ram[6671]  = 252;
  ram[6672]  = 255;
  ram[6673]  = 255;
  ram[6674]  = 255;
  ram[6675]  = 255;
  ram[6676]  = 255;
  ram[6677]  = 255;
  ram[6678]  = 254;
  ram[6679]  = 254;
  ram[6680]  = 255;
  ram[6681]  = 255;
  ram[6682]  = 255;
  ram[6683]  = 255;
  ram[6684]  = 252;
  ram[6685]  = 255;
  ram[6686]  = 255;
  ram[6687]  = 255;
  ram[6688]  = 255;
  ram[6689]  = 255;
  ram[6690]  = 255;
  ram[6691]  = 255;
  ram[6692]  = 254;
  ram[6693]  = 254;
  ram[6694]  = 253;
  ram[6695]  = 250;
  ram[6696]  = 255;
  ram[6697]  = 255;
  ram[6698]  = 255;
  ram[6699]  = 255;
  ram[6700]  = 255;
  ram[6701]  = 255;
  ram[6702]  = 247;
  ram[6703]  = 252;
  ram[6704]  = 251;
  ram[6705]  = 255;
  ram[6706]  = 255;
  ram[6707]  = 255;
  ram[6708]  = 254;
  ram[6709]  = 253;
  ram[6710]  = 250;
  ram[6711]  = 255;
  ram[6712]  = 255;
  ram[6713]  = 255;
  ram[6714]  = 254;
  ram[6715]  = 255;
  ram[6716]  = 255;
  ram[6717]  = 255;
  ram[6718]  = 255;
  ram[6719]  = 255;
  ram[6720]  = 255;
  ram[6721]  = 255;
  ram[6722]  = 253;
  ram[6723]  = 254;
  ram[6724]  = 254;
  ram[6725]  = 255;
  ram[6726]  = 255;
  ram[6727]  = 255;
  ram[6728]  = 253;
  ram[6729]  = 249;
  ram[6730]  = 255;
  ram[6731]  = 255;
  ram[6732]  = 249;
  ram[6733]  = 253;
  ram[6734]  = 255;
  ram[6735]  = 255;
  ram[6736]  = 255;
  ram[6737]  = 255;
  ram[6738]  = 254;
  ram[6739]  = 255;
  ram[6740]  = 255;
  ram[6741]  = 255;
  ram[6742]  = 255;
  ram[6743]  = 251;
  ram[6744]  = 252;
  ram[6745]  = 255;
  ram[6746]  = 255;
  ram[6747]  = 255;
  ram[6748]  = 255;
  ram[6749]  = 255;
  ram[6750]  = 253;
  ram[6751]  = 253;
  ram[6752]  = 255;
  ram[6753]  = 255;
  ram[6754]  = 255;
  ram[6755]  = 255;
  ram[6756]  = 253;
  ram[6757]  = 255;
  ram[6758]  = 255;
  ram[6759]  = 255;
  ram[6760]  = 255;
  ram[6761]  = 255;
  ram[6762]  = 252;
  ram[6763]  = 250;
  ram[6764]  = 251;
  ram[6765]  = 253;
  ram[6766]  = 255;
  ram[6767]  = 255;
  ram[6768]  = 255;
  ram[6769]  = 250;
  ram[6770]  = 255;
  ram[6771]  = 255;
  ram[6772]  = 255;
  ram[6773]  = 255;
  ram[6774]  = 253;
  ram[6775]  = 255;
  ram[6776]  = 255;
  ram[6777]  = 253;
  ram[6778]  = 255;
  ram[6779]  = 255;
  ram[6780]  = 253;
  ram[6781]  = 255;
  ram[6782]  = 255;
  ram[6783]  = 253;
  ram[6784]  = 251;
  ram[6785]  = 255;
  ram[6786]  = 255;
  ram[6787]  = 255;
  ram[6788]  = 255;
  ram[6789]  = 255;
  ram[6790]  = 255;
  ram[6791]  = 255;
  ram[6792]  = 255;
  ram[6793]  = 255;
  ram[6794]  = 255;
  ram[6795]  = 255;
  ram[6796]  = 236;
  ram[6797]  = 211;
  ram[6798]  = 243;
  ram[6799]  = 255;
  ram[6800]  = 253;
  ram[6801]  = 235;
  ram[6802]  = 209;
  ram[6803]  = 242;
  ram[6804]  = 255;
  ram[6805]  = 254;
  ram[6806]  = 252;
  ram[6807]  = 255;
  ram[6808]  = 255;
  ram[6809]  = 255;
  ram[6810]  = 255;
  ram[6811]  = 255;
  ram[6812]  = 255;
  ram[6813]  = 255;
  ram[6814]  = 254;
  ram[6815]  = 252;
  ram[6816]  = 254;
  ram[6817]  = 254;
  ram[6818]  = 253;
  ram[6819]  = 253;
  ram[6820]  = 255;
  ram[6821]  = 255;
  ram[6822]  = 255;
  ram[6823]  = 255;
  ram[6824]  = 253;
  ram[6825]  = 253;
  ram[6826]  = 253;
  ram[6827]  = 253;
  ram[6828]  = 252;
  ram[6829]  = 255;
  ram[6830]  = 255;
  ram[6831]  = 255;
  ram[6832]  = 253;
  ram[6833]  = 252;
  ram[6834]  = 254;
  ram[6835]  = 253;
  ram[6836]  = 254;
  ram[6837]  = 251;
  ram[6838]  = 252;
  ram[6839]  = 254;
  ram[6840]  = 252;
  ram[6841]  = 251;
  ram[6842]  = 254;
  ram[6843]  = 254;
  ram[6844]  = 252;
  ram[6845]  = 252;
  ram[6846]  = 252;
  ram[6847]  = 254;
  ram[6848]  = 255;
  ram[6849]  = 252;
  ram[6850]  = 254;
  ram[6851]  = 253;
  ram[6852]  = 255;
  ram[6853]  = 255;
  ram[6854]  = 255;
  ram[6855]  = 255;
  ram[6856]  = 253;
  ram[6857]  = 254;
  ram[6858]  = 253;
  ram[6859]  = 253;
  ram[6860]  = 254;
  ram[6861]  = 252;
  ram[6862]  = 253;
  ram[6863]  = 253;
  ram[6864]  = 253;
  ram[6865]  = 252;
  ram[6866]  = 254;
  ram[6867]  = 252;
  ram[6868]  = 253;
  ram[6869]  = 252;
  ram[6870]  = 254;
  ram[6871]  = 252;
  ram[6872]  = 252;
  ram[6873]  = 253;
  ram[6874]  = 253;
  ram[6875]  = 253;
  ram[6876]  = 254;
  ram[6877]  = 254;
  ram[6878]  = 254;
  ram[6879]  = 254;
  ram[6880]  = 255;
  ram[6881]  = 255;
  ram[6882]  = 255;
  ram[6883]  = 255;
  ram[6884]  = 255;
  ram[6885]  = 253;
  ram[6886]  = 254;
  ram[6887]  = 253;
  ram[6888]  = 253;
  ram[6889]  = 252;
  ram[6890]  = 254;
  ram[6891]  = 253;
  ram[6892]  = 253;
  ram[6893]  = 255;
  ram[6894]  = 254;
  ram[6895]  = 252;
  ram[6896]  = 252;
  ram[6897]  = 254;
  ram[6898]  = 254;
  ram[6899]  = 253;
  ram[6900]  = 252;
  ram[6901]  = 253;
  ram[6902]  = 251;
  ram[6903]  = 253;
  ram[6904]  = 251;
  ram[6905]  = 253;
  ram[6906]  = 252;
  ram[6907]  = 254;
  ram[6908]  = 253;
  ram[6909]  = 252;
  ram[6910]  = 251;
  ram[6911]  = 253;
  ram[6912]  = 252;
  ram[6913]  = 253;
  ram[6914]  = 255;
  ram[6915]  = 255;
  ram[6916]  = 253;
  ram[6917]  = 251;
  ram[6918]  = 253;
  ram[6919]  = 253;
  ram[6920]  = 253;
  ram[6921]  = 253;
  ram[6922]  = 254;
  ram[6923]  = 253;
  ram[6924]  = 253;
  ram[6925]  = 252;
  ram[6926]  = 254;
  ram[6927]  = 253;
  ram[6928]  = 252;
  ram[6929]  = 252;
  ram[6930]  = 253;
  ram[6931]  = 254;
  ram[6932]  = 252;
  ram[6933]  = 254;
  ram[6934]  = 255;
  ram[6935]  = 255;
  ram[6936]  = 255;
  ram[6937]  = 255;
  ram[6938]  = 253;
  ram[6939]  = 252;
  ram[6940]  = 251;
  ram[6941]  = 253;
  ram[6942]  = 253;
  ram[6943]  = 252;
  ram[6944]  = 253;
  ram[6945]  = 251;
  ram[6946]  = 253;
  ram[6947]  = 252;
  ram[6948]  = 254;
  ram[6949]  = 252;
  ram[6950]  = 253;
  ram[6951]  = 255;
  ram[6952]  = 255;
  ram[6953]  = 255;
  ram[6954]  = 255;
  ram[6955]  = 255;
  ram[6956]  = 254;
  ram[6957]  = 253;
  ram[6958]  = 252;
  ram[6959]  = 252;
  ram[6960]  = 253;
  ram[6961]  = 253;
  ram[6962]  = 254;
  ram[6963]  = 252;
  ram[6964]  = 254;
  ram[6965]  = 252;
  ram[6966]  = 252;
  ram[6967]  = 253;
  ram[6968]  = 253;
  ram[6969]  = 251;
  ram[6970]  = 251;
  ram[6971]  = 253;
  ram[6972]  = 253;
  ram[6973]  = 252;
  ram[6974]  = 253;
  ram[6975]  = 253;
  ram[6976]  = 252;
  ram[6977]  = 252;
  ram[6978]  = 254;
  ram[6979]  = 252;
  ram[6980]  = 252;
  ram[6981]  = 255;
  ram[6982]  = 255;
  ram[6983]  = 252;
  ram[6984]  = 254;
  ram[6985]  = 250;
  ram[6986]  = 250;
  ram[6987]  = 251;
  ram[6988]  = 254;
  ram[6989]  = 255;
  ram[6990]  = 255;
  ram[6991]  = 255;
  ram[6992]  = 255;
  ram[6993]  = 255;
  ram[6994]  = 255;
  ram[6995]  = 255;
  ram[6996]  = 236;
  ram[6997]  = 211;
  ram[6998]  = 243;
  ram[6999]  = 255;
  ram[7000]  = 253;
  ram[7001]  = 235;
  ram[7002]  = 209;
  ram[7003]  = 242;
  ram[7004]  = 255;
  ram[7005]  = 254;
  ram[7006]  = 252;
  ram[7007]  = 255;
  ram[7008]  = 255;
  ram[7009]  = 255;
  ram[7010]  = 255;
  ram[7011]  = 255;
  ram[7012]  = 255;
  ram[7013]  = 255;
  ram[7014]  = 255;
  ram[7015]  = 254;
  ram[7016]  = 255;
  ram[7017]  = 255;
  ram[7018]  = 255;
  ram[7019]  = 255;
  ram[7020]  = 255;
  ram[7021]  = 255;
  ram[7022]  = 255;
  ram[7023]  = 255;
  ram[7024]  = 255;
  ram[7025]  = 255;
  ram[7026]  = 254;
  ram[7027]  = 254;
  ram[7028]  = 254;
  ram[7029]  = 255;
  ram[7030]  = 255;
  ram[7031]  = 255;
  ram[7032]  = 255;
  ram[7033]  = 254;
  ram[7034]  = 255;
  ram[7035]  = 255;
  ram[7036]  = 255;
  ram[7037]  = 254;
  ram[7038]  = 254;
  ram[7039]  = 254;
  ram[7040]  = 254;
  ram[7041]  = 254;
  ram[7042]  = 255;
  ram[7043]  = 255;
  ram[7044]  = 254;
  ram[7045]  = 254;
  ram[7046]  = 254;
  ram[7047]  = 255;
  ram[7048]  = 255;
  ram[7049]  = 254;
  ram[7050]  = 254;
  ram[7051]  = 254;
  ram[7052]  = 255;
  ram[7053]  = 255;
  ram[7054]  = 255;
  ram[7055]  = 255;
  ram[7056]  = 254;
  ram[7057]  = 254;
  ram[7058]  = 254;
  ram[7059]  = 254;
  ram[7060]  = 255;
  ram[7061]  = 254;
  ram[7062]  = 254;
  ram[7063]  = 254;
  ram[7064]  = 255;
  ram[7065]  = 254;
  ram[7066]  = 254;
  ram[7067]  = 254;
  ram[7068]  = 254;
  ram[7069]  = 254;
  ram[7070]  = 254;
  ram[7071]  = 255;
  ram[7072]  = 254;
  ram[7073]  = 254;
  ram[7074]  = 255;
  ram[7075]  = 255;
  ram[7076]  = 255;
  ram[7077]  = 255;
  ram[7078]  = 254;
  ram[7079]  = 255;
  ram[7080]  = 255;
  ram[7081]  = 255;
  ram[7082]  = 255;
  ram[7083]  = 255;
  ram[7084]  = 255;
  ram[7085]  = 254;
  ram[7086]  = 255;
  ram[7087]  = 255;
  ram[7088]  = 254;
  ram[7089]  = 255;
  ram[7090]  = 254;
  ram[7091]  = 254;
  ram[7092]  = 254;
  ram[7093]  = 255;
  ram[7094]  = 255;
  ram[7095]  = 255;
  ram[7096]  = 255;
  ram[7097]  = 255;
  ram[7098]  = 255;
  ram[7099]  = 254;
  ram[7100]  = 255;
  ram[7101]  = 254;
  ram[7102]  = 254;
  ram[7103]  = 255;
  ram[7104]  = 255;
  ram[7105]  = 255;
  ram[7106]  = 254;
  ram[7107]  = 255;
  ram[7108]  = 255;
  ram[7109]  = 255;
  ram[7110]  = 255;
  ram[7111]  = 254;
  ram[7112]  = 254;
  ram[7113]  = 254;
  ram[7114]  = 255;
  ram[7115]  = 255;
  ram[7116]  = 255;
  ram[7117]  = 254;
  ram[7118]  = 254;
  ram[7119]  = 255;
  ram[7120]  = 255;
  ram[7121]  = 255;
  ram[7122]  = 255;
  ram[7123]  = 254;
  ram[7124]  = 254;
  ram[7125]  = 254;
  ram[7126]  = 255;
  ram[7127]  = 254;
  ram[7128]  = 254;
  ram[7129]  = 254;
  ram[7130]  = 254;
  ram[7131]  = 255;
  ram[7132]  = 254;
  ram[7133]  = 255;
  ram[7134]  = 255;
  ram[7135]  = 255;
  ram[7136]  = 255;
  ram[7137]  = 255;
  ram[7138]  = 255;
  ram[7139]  = 255;
  ram[7140]  = 254;
  ram[7141]  = 254;
  ram[7142]  = 254;
  ram[7143]  = 254;
  ram[7144]  = 254;
  ram[7145]  = 255;
  ram[7146]  = 254;
  ram[7147]  = 254;
  ram[7148]  = 255;
  ram[7149]  = 254;
  ram[7150]  = 255;
  ram[7151]  = 255;
  ram[7152]  = 255;
  ram[7153]  = 255;
  ram[7154]  = 255;
  ram[7155]  = 255;
  ram[7156]  = 255;
  ram[7157]  = 254;
  ram[7158]  = 254;
  ram[7159]  = 254;
  ram[7160]  = 254;
  ram[7161]  = 255;
  ram[7162]  = 254;
  ram[7163]  = 255;
  ram[7164]  = 255;
  ram[7165]  = 254;
  ram[7166]  = 255;
  ram[7167]  = 255;
  ram[7168]  = 255;
  ram[7169]  = 255;
  ram[7170]  = 254;
  ram[7171]  = 254;
  ram[7172]  = 255;
  ram[7173]  = 254;
  ram[7174]  = 254;
  ram[7175]  = 255;
  ram[7176]  = 255;
  ram[7177]  = 254;
  ram[7178]  = 255;
  ram[7179]  = 254;
  ram[7180]  = 254;
  ram[7181]  = 255;
  ram[7182]  = 255;
  ram[7183]  = 255;
  ram[7184]  = 254;
  ram[7185]  = 255;
  ram[7186]  = 254;
  ram[7187]  = 255;
  ram[7188]  = 255;
  ram[7189]  = 255;
  ram[7190]  = 255;
  ram[7191]  = 255;
  ram[7192]  = 255;
  ram[7193]  = 255;
  ram[7194]  = 255;
  ram[7195]  = 255;
  ram[7196]  = 236;
  ram[7197]  = 211;
  ram[7198]  = 243;
  ram[7199]  = 255;
  ram[7200]  = 253;
  ram[7201]  = 235;
  ram[7202]  = 209;
  ram[7203]  = 242;
  ram[7204]  = 255;
  ram[7205]  = 254;
  ram[7206]  = 252;
  ram[7207]  = 255;
  ram[7208]  = 255;
  ram[7209]  = 255;
  ram[7210]  = 255;
  ram[7211]  = 255;
  ram[7212]  = 255;
  ram[7213]  = 255;
  ram[7214]  = 255;
  ram[7215]  = 255;
  ram[7216]  = 255;
  ram[7217]  = 255;
  ram[7218]  = 255;
  ram[7219]  = 255;
  ram[7220]  = 255;
  ram[7221]  = 255;
  ram[7222]  = 255;
  ram[7223]  = 255;
  ram[7224]  = 255;
  ram[7225]  = 255;
  ram[7226]  = 255;
  ram[7227]  = 255;
  ram[7228]  = 255;
  ram[7229]  = 255;
  ram[7230]  = 255;
  ram[7231]  = 255;
  ram[7232]  = 255;
  ram[7233]  = 255;
  ram[7234]  = 255;
  ram[7235]  = 255;
  ram[7236]  = 255;
  ram[7237]  = 255;
  ram[7238]  = 255;
  ram[7239]  = 255;
  ram[7240]  = 255;
  ram[7241]  = 255;
  ram[7242]  = 255;
  ram[7243]  = 255;
  ram[7244]  = 255;
  ram[7245]  = 255;
  ram[7246]  = 255;
  ram[7247]  = 255;
  ram[7248]  = 255;
  ram[7249]  = 255;
  ram[7250]  = 255;
  ram[7251]  = 255;
  ram[7252]  = 255;
  ram[7253]  = 255;
  ram[7254]  = 255;
  ram[7255]  = 255;
  ram[7256]  = 255;
  ram[7257]  = 255;
  ram[7258]  = 255;
  ram[7259]  = 255;
  ram[7260]  = 255;
  ram[7261]  = 255;
  ram[7262]  = 255;
  ram[7263]  = 255;
  ram[7264]  = 255;
  ram[7265]  = 255;
  ram[7266]  = 255;
  ram[7267]  = 255;
  ram[7268]  = 255;
  ram[7269]  = 255;
  ram[7270]  = 255;
  ram[7271]  = 255;
  ram[7272]  = 255;
  ram[7273]  = 255;
  ram[7274]  = 255;
  ram[7275]  = 255;
  ram[7276]  = 255;
  ram[7277]  = 255;
  ram[7278]  = 255;
  ram[7279]  = 255;
  ram[7280]  = 255;
  ram[7281]  = 255;
  ram[7282]  = 255;
  ram[7283]  = 255;
  ram[7284]  = 255;
  ram[7285]  = 255;
  ram[7286]  = 255;
  ram[7287]  = 255;
  ram[7288]  = 255;
  ram[7289]  = 255;
  ram[7290]  = 255;
  ram[7291]  = 255;
  ram[7292]  = 255;
  ram[7293]  = 255;
  ram[7294]  = 255;
  ram[7295]  = 255;
  ram[7296]  = 255;
  ram[7297]  = 255;
  ram[7298]  = 255;
  ram[7299]  = 255;
  ram[7300]  = 255;
  ram[7301]  = 255;
  ram[7302]  = 255;
  ram[7303]  = 255;
  ram[7304]  = 255;
  ram[7305]  = 255;
  ram[7306]  = 255;
  ram[7307]  = 255;
  ram[7308]  = 255;
  ram[7309]  = 255;
  ram[7310]  = 255;
  ram[7311]  = 255;
  ram[7312]  = 255;
  ram[7313]  = 255;
  ram[7314]  = 255;
  ram[7315]  = 255;
  ram[7316]  = 255;
  ram[7317]  = 255;
  ram[7318]  = 255;
  ram[7319]  = 255;
  ram[7320]  = 255;
  ram[7321]  = 255;
  ram[7322]  = 255;
  ram[7323]  = 255;
  ram[7324]  = 255;
  ram[7325]  = 255;
  ram[7326]  = 255;
  ram[7327]  = 255;
  ram[7328]  = 255;
  ram[7329]  = 255;
  ram[7330]  = 255;
  ram[7331]  = 255;
  ram[7332]  = 255;
  ram[7333]  = 255;
  ram[7334]  = 255;
  ram[7335]  = 255;
  ram[7336]  = 255;
  ram[7337]  = 255;
  ram[7338]  = 255;
  ram[7339]  = 255;
  ram[7340]  = 255;
  ram[7341]  = 255;
  ram[7342]  = 255;
  ram[7343]  = 255;
  ram[7344]  = 255;
  ram[7345]  = 255;
  ram[7346]  = 255;
  ram[7347]  = 255;
  ram[7348]  = 255;
  ram[7349]  = 255;
  ram[7350]  = 255;
  ram[7351]  = 255;
  ram[7352]  = 255;
  ram[7353]  = 255;
  ram[7354]  = 255;
  ram[7355]  = 255;
  ram[7356]  = 255;
  ram[7357]  = 255;
  ram[7358]  = 255;
  ram[7359]  = 255;
  ram[7360]  = 255;
  ram[7361]  = 255;
  ram[7362]  = 255;
  ram[7363]  = 255;
  ram[7364]  = 255;
  ram[7365]  = 255;
  ram[7366]  = 255;
  ram[7367]  = 255;
  ram[7368]  = 255;
  ram[7369]  = 255;
  ram[7370]  = 255;
  ram[7371]  = 255;
  ram[7372]  = 255;
  ram[7373]  = 255;
  ram[7374]  = 255;
  ram[7375]  = 255;
  ram[7376]  = 255;
  ram[7377]  = 255;
  ram[7378]  = 255;
  ram[7379]  = 255;
  ram[7380]  = 255;
  ram[7381]  = 255;
  ram[7382]  = 255;
  ram[7383]  = 255;
  ram[7384]  = 255;
  ram[7385]  = 255;
  ram[7386]  = 255;
  ram[7387]  = 255;
  ram[7388]  = 255;
  ram[7389]  = 255;
  ram[7390]  = 255;
  ram[7391]  = 255;
  ram[7392]  = 255;
  ram[7393]  = 255;
  ram[7394]  = 255;
  ram[7395]  = 255;
  ram[7396]  = 236;
  ram[7397]  = 211;
  ram[7398]  = 243;
  ram[7399]  = 255;
  ram[7400]  = 252;
  ram[7401]  = 235;
  ram[7402]  = 209;
  ram[7403]  = 242;
  ram[7404]  = 255;
  ram[7405]  = 254;
  ram[7406]  = 252;
  ram[7407]  = 255;
  ram[7408]  = 255;
  ram[7409]  = 255;
  ram[7410]  = 255;
  ram[7411]  = 255;
  ram[7412]  = 255;
  ram[7413]  = 255;
  ram[7414]  = 255;
  ram[7415]  = 255;
  ram[7416]  = 255;
  ram[7417]  = 255;
  ram[7418]  = 255;
  ram[7419]  = 255;
  ram[7420]  = 255;
  ram[7421]  = 255;
  ram[7422]  = 255;
  ram[7423]  = 255;
  ram[7424]  = 255;
  ram[7425]  = 255;
  ram[7426]  = 255;
  ram[7427]  = 255;
  ram[7428]  = 255;
  ram[7429]  = 255;
  ram[7430]  = 255;
  ram[7431]  = 255;
  ram[7432]  = 255;
  ram[7433]  = 255;
  ram[7434]  = 255;
  ram[7435]  = 255;
  ram[7436]  = 255;
  ram[7437]  = 255;
  ram[7438]  = 255;
  ram[7439]  = 255;
  ram[7440]  = 255;
  ram[7441]  = 255;
  ram[7442]  = 255;
  ram[7443]  = 255;
  ram[7444]  = 255;
  ram[7445]  = 255;
  ram[7446]  = 255;
  ram[7447]  = 255;
  ram[7448]  = 255;
  ram[7449]  = 255;
  ram[7450]  = 255;
  ram[7451]  = 255;
  ram[7452]  = 255;
  ram[7453]  = 255;
  ram[7454]  = 255;
  ram[7455]  = 255;
  ram[7456]  = 255;
  ram[7457]  = 255;
  ram[7458]  = 255;
  ram[7459]  = 255;
  ram[7460]  = 255;
  ram[7461]  = 255;
  ram[7462]  = 255;
  ram[7463]  = 255;
  ram[7464]  = 255;
  ram[7465]  = 255;
  ram[7466]  = 255;
  ram[7467]  = 255;
  ram[7468]  = 255;
  ram[7469]  = 255;
  ram[7470]  = 255;
  ram[7471]  = 255;
  ram[7472]  = 255;
  ram[7473]  = 255;
  ram[7474]  = 255;
  ram[7475]  = 255;
  ram[7476]  = 255;
  ram[7477]  = 255;
  ram[7478]  = 255;
  ram[7479]  = 255;
  ram[7480]  = 255;
  ram[7481]  = 255;
  ram[7482]  = 255;
  ram[7483]  = 255;
  ram[7484]  = 255;
  ram[7485]  = 255;
  ram[7486]  = 255;
  ram[7487]  = 255;
  ram[7488]  = 255;
  ram[7489]  = 255;
  ram[7490]  = 255;
  ram[7491]  = 255;
  ram[7492]  = 255;
  ram[7493]  = 255;
  ram[7494]  = 255;
  ram[7495]  = 255;
  ram[7496]  = 255;
  ram[7497]  = 255;
  ram[7498]  = 255;
  ram[7499]  = 255;
  ram[7500]  = 255;
  ram[7501]  = 255;
  ram[7502]  = 255;
  ram[7503]  = 255;
  ram[7504]  = 255;
  ram[7505]  = 255;
  ram[7506]  = 255;
  ram[7507]  = 255;
  ram[7508]  = 255;
  ram[7509]  = 255;
  ram[7510]  = 255;
  ram[7511]  = 255;
  ram[7512]  = 255;
  ram[7513]  = 255;
  ram[7514]  = 255;
  ram[7515]  = 255;
  ram[7516]  = 255;
  ram[7517]  = 255;
  ram[7518]  = 255;
  ram[7519]  = 255;
  ram[7520]  = 255;
  ram[7521]  = 255;
  ram[7522]  = 255;
  ram[7523]  = 255;
  ram[7524]  = 255;
  ram[7525]  = 255;
  ram[7526]  = 255;
  ram[7527]  = 255;
  ram[7528]  = 255;
  ram[7529]  = 255;
  ram[7530]  = 255;
  ram[7531]  = 255;
  ram[7532]  = 255;
  ram[7533]  = 255;
  ram[7534]  = 255;
  ram[7535]  = 255;
  ram[7536]  = 255;
  ram[7537]  = 255;
  ram[7538]  = 255;
  ram[7539]  = 255;
  ram[7540]  = 255;
  ram[7541]  = 255;
  ram[7542]  = 255;
  ram[7543]  = 255;
  ram[7544]  = 255;
  ram[7545]  = 255;
  ram[7546]  = 255;
  ram[7547]  = 255;
  ram[7548]  = 255;
  ram[7549]  = 255;
  ram[7550]  = 255;
  ram[7551]  = 255;
  ram[7552]  = 255;
  ram[7553]  = 255;
  ram[7554]  = 255;
  ram[7555]  = 255;
  ram[7556]  = 255;
  ram[7557]  = 255;
  ram[7558]  = 255;
  ram[7559]  = 255;
  ram[7560]  = 255;
  ram[7561]  = 255;
  ram[7562]  = 255;
  ram[7563]  = 255;
  ram[7564]  = 255;
  ram[7565]  = 255;
  ram[7566]  = 255;
  ram[7567]  = 255;
  ram[7568]  = 255;
  ram[7569]  = 255;
  ram[7570]  = 255;
  ram[7571]  = 255;
  ram[7572]  = 255;
  ram[7573]  = 255;
  ram[7574]  = 255;
  ram[7575]  = 255;
  ram[7576]  = 255;
  ram[7577]  = 255;
  ram[7578]  = 255;
  ram[7579]  = 255;
  ram[7580]  = 255;
  ram[7581]  = 255;
  ram[7582]  = 255;
  ram[7583]  = 255;
  ram[7584]  = 255;
  ram[7585]  = 255;
  ram[7586]  = 255;
  ram[7587]  = 255;
  ram[7588]  = 255;
  ram[7589]  = 255;
  ram[7590]  = 255;
  ram[7591]  = 255;
  ram[7592]  = 255;
  ram[7593]  = 255;
  ram[7594]  = 255;
  ram[7595]  = 255;
  ram[7596]  = 236;
  ram[7597]  = 211;
  ram[7598]  = 243;
  ram[7599]  = 255;
  ram[7600]  = 255;
  ram[7601]  = 234;
  ram[7602]  = 205;
  ram[7603]  = 242;
  ram[7604]  = 255;
  ram[7605]  = 254;
  ram[7606]  = 251;
  ram[7607]  = 255;
  ram[7608]  = 255;
  ram[7609]  = 255;
  ram[7610]  = 255;
  ram[7611]  = 255;
  ram[7612]  = 255;
  ram[7613]  = 255;
  ram[7614]  = 255;
  ram[7615]  = 255;
  ram[7616]  = 255;
  ram[7617]  = 255;
  ram[7618]  = 255;
  ram[7619]  = 255;
  ram[7620]  = 255;
  ram[7621]  = 255;
  ram[7622]  = 255;
  ram[7623]  = 255;
  ram[7624]  = 255;
  ram[7625]  = 255;
  ram[7626]  = 255;
  ram[7627]  = 255;
  ram[7628]  = 255;
  ram[7629]  = 255;
  ram[7630]  = 255;
  ram[7631]  = 255;
  ram[7632]  = 255;
  ram[7633]  = 255;
  ram[7634]  = 255;
  ram[7635]  = 255;
  ram[7636]  = 255;
  ram[7637]  = 255;
  ram[7638]  = 255;
  ram[7639]  = 255;
  ram[7640]  = 255;
  ram[7641]  = 255;
  ram[7642]  = 255;
  ram[7643]  = 255;
  ram[7644]  = 255;
  ram[7645]  = 255;
  ram[7646]  = 255;
  ram[7647]  = 255;
  ram[7648]  = 255;
  ram[7649]  = 255;
  ram[7650]  = 255;
  ram[7651]  = 255;
  ram[7652]  = 255;
  ram[7653]  = 255;
  ram[7654]  = 255;
  ram[7655]  = 255;
  ram[7656]  = 255;
  ram[7657]  = 255;
  ram[7658]  = 255;
  ram[7659]  = 255;
  ram[7660]  = 255;
  ram[7661]  = 255;
  ram[7662]  = 255;
  ram[7663]  = 255;
  ram[7664]  = 255;
  ram[7665]  = 255;
  ram[7666]  = 255;
  ram[7667]  = 255;
  ram[7668]  = 255;
  ram[7669]  = 255;
  ram[7670]  = 255;
  ram[7671]  = 255;
  ram[7672]  = 255;
  ram[7673]  = 255;
  ram[7674]  = 255;
  ram[7675]  = 255;
  ram[7676]  = 255;
  ram[7677]  = 255;
  ram[7678]  = 255;
  ram[7679]  = 255;
  ram[7680]  = 255;
  ram[7681]  = 255;
  ram[7682]  = 255;
  ram[7683]  = 255;
  ram[7684]  = 255;
  ram[7685]  = 255;
  ram[7686]  = 255;
  ram[7687]  = 255;
  ram[7688]  = 255;
  ram[7689]  = 255;
  ram[7690]  = 255;
  ram[7691]  = 255;
  ram[7692]  = 255;
  ram[7693]  = 255;
  ram[7694]  = 255;
  ram[7695]  = 255;
  ram[7696]  = 255;
  ram[7697]  = 255;
  ram[7698]  = 255;
  ram[7699]  = 255;
  ram[7700]  = 255;
  ram[7701]  = 255;
  ram[7702]  = 255;
  ram[7703]  = 255;
  ram[7704]  = 255;
  ram[7705]  = 255;
  ram[7706]  = 255;
  ram[7707]  = 255;
  ram[7708]  = 255;
  ram[7709]  = 255;
  ram[7710]  = 255;
  ram[7711]  = 255;
  ram[7712]  = 255;
  ram[7713]  = 255;
  ram[7714]  = 255;
  ram[7715]  = 255;
  ram[7716]  = 255;
  ram[7717]  = 255;
  ram[7718]  = 255;
  ram[7719]  = 255;
  ram[7720]  = 255;
  ram[7721]  = 255;
  ram[7722]  = 255;
  ram[7723]  = 255;
  ram[7724]  = 255;
  ram[7725]  = 255;
  ram[7726]  = 255;
  ram[7727]  = 255;
  ram[7728]  = 255;
  ram[7729]  = 255;
  ram[7730]  = 255;
  ram[7731]  = 255;
  ram[7732]  = 255;
  ram[7733]  = 255;
  ram[7734]  = 255;
  ram[7735]  = 255;
  ram[7736]  = 255;
  ram[7737]  = 255;
  ram[7738]  = 255;
  ram[7739]  = 255;
  ram[7740]  = 255;
  ram[7741]  = 255;
  ram[7742]  = 255;
  ram[7743]  = 255;
  ram[7744]  = 255;
  ram[7745]  = 255;
  ram[7746]  = 255;
  ram[7747]  = 255;
  ram[7748]  = 255;
  ram[7749]  = 255;
  ram[7750]  = 255;
  ram[7751]  = 255;
  ram[7752]  = 255;
  ram[7753]  = 255;
  ram[7754]  = 255;
  ram[7755]  = 255;
  ram[7756]  = 255;
  ram[7757]  = 255;
  ram[7758]  = 255;
  ram[7759]  = 255;
  ram[7760]  = 255;
  ram[7761]  = 255;
  ram[7762]  = 255;
  ram[7763]  = 255;
  ram[7764]  = 255;
  ram[7765]  = 255;
  ram[7766]  = 255;
  ram[7767]  = 255;
  ram[7768]  = 255;
  ram[7769]  = 255;
  ram[7770]  = 255;
  ram[7771]  = 255;
  ram[7772]  = 255;
  ram[7773]  = 255;
  ram[7774]  = 255;
  ram[7775]  = 255;
  ram[7776]  = 255;
  ram[7777]  = 255;
  ram[7778]  = 255;
  ram[7779]  = 255;
  ram[7780]  = 255;
  ram[7781]  = 255;
  ram[7782]  = 255;
  ram[7783]  = 255;
  ram[7784]  = 255;
  ram[7785]  = 255;
  ram[7786]  = 255;
  ram[7787]  = 255;
  ram[7788]  = 255;
  ram[7789]  = 255;
  ram[7790]  = 255;
  ram[7791]  = 255;
  ram[7792]  = 255;
  ram[7793]  = 255;
  ram[7794]  = 255;
  ram[7795]  = 255;
  ram[7796]  = 236;
  ram[7797]  = 212;
  ram[7798]  = 243;
  ram[7799]  = 255;
  ram[7800]  = 255;
  ram[7801]  = 232;
  ram[7802]  = 204;
  ram[7803]  = 243;
  ram[7804]  = 255;
  ram[7805]  = 254;
  ram[7806]  = 251;
  ram[7807]  = 255;
  ram[7808]  = 255;
  ram[7809]  = 255;
  ram[7810]  = 255;
  ram[7811]  = 255;
  ram[7812]  = 255;
  ram[7813]  = 255;
  ram[7814]  = 255;
  ram[7815]  = 255;
  ram[7816]  = 255;
  ram[7817]  = 255;
  ram[7818]  = 255;
  ram[7819]  = 255;
  ram[7820]  = 255;
  ram[7821]  = 255;
  ram[7822]  = 255;
  ram[7823]  = 255;
  ram[7824]  = 255;
  ram[7825]  = 255;
  ram[7826]  = 255;
  ram[7827]  = 255;
  ram[7828]  = 255;
  ram[7829]  = 255;
  ram[7830]  = 255;
  ram[7831]  = 255;
  ram[7832]  = 255;
  ram[7833]  = 255;
  ram[7834]  = 255;
  ram[7835]  = 255;
  ram[7836]  = 255;
  ram[7837]  = 255;
  ram[7838]  = 255;
  ram[7839]  = 255;
  ram[7840]  = 255;
  ram[7841]  = 255;
  ram[7842]  = 255;
  ram[7843]  = 255;
  ram[7844]  = 255;
  ram[7845]  = 255;
  ram[7846]  = 255;
  ram[7847]  = 255;
  ram[7848]  = 255;
  ram[7849]  = 255;
  ram[7850]  = 255;
  ram[7851]  = 255;
  ram[7852]  = 255;
  ram[7853]  = 255;
  ram[7854]  = 255;
  ram[7855]  = 255;
  ram[7856]  = 255;
  ram[7857]  = 255;
  ram[7858]  = 255;
  ram[7859]  = 255;
  ram[7860]  = 255;
  ram[7861]  = 255;
  ram[7862]  = 255;
  ram[7863]  = 255;
  ram[7864]  = 255;
  ram[7865]  = 255;
  ram[7866]  = 255;
  ram[7867]  = 255;
  ram[7868]  = 255;
  ram[7869]  = 255;
  ram[7870]  = 255;
  ram[7871]  = 255;
  ram[7872]  = 255;
  ram[7873]  = 255;
  ram[7874]  = 255;
  ram[7875]  = 255;
  ram[7876]  = 255;
  ram[7877]  = 255;
  ram[7878]  = 255;
  ram[7879]  = 255;
  ram[7880]  = 255;
  ram[7881]  = 255;
  ram[7882]  = 255;
  ram[7883]  = 255;
  ram[7884]  = 255;
  ram[7885]  = 255;
  ram[7886]  = 255;
  ram[7887]  = 255;
  ram[7888]  = 255;
  ram[7889]  = 255;
  ram[7890]  = 255;
  ram[7891]  = 255;
  ram[7892]  = 255;
  ram[7893]  = 255;
  ram[7894]  = 255;
  ram[7895]  = 255;
  ram[7896]  = 255;
  ram[7897]  = 255;
  ram[7898]  = 255;
  ram[7899]  = 255;
  ram[7900]  = 255;
  ram[7901]  = 255;
  ram[7902]  = 255;
  ram[7903]  = 255;
  ram[7904]  = 255;
  ram[7905]  = 255;
  ram[7906]  = 255;
  ram[7907]  = 255;
  ram[7908]  = 255;
  ram[7909]  = 255;
  ram[7910]  = 255;
  ram[7911]  = 255;
  ram[7912]  = 255;
  ram[7913]  = 255;
  ram[7914]  = 255;
  ram[7915]  = 255;
  ram[7916]  = 255;
  ram[7917]  = 255;
  ram[7918]  = 255;
  ram[7919]  = 255;
  ram[7920]  = 255;
  ram[7921]  = 255;
  ram[7922]  = 255;
  ram[7923]  = 255;
  ram[7924]  = 255;
  ram[7925]  = 255;
  ram[7926]  = 255;
  ram[7927]  = 255;
  ram[7928]  = 255;
  ram[7929]  = 255;
  ram[7930]  = 255;
  ram[7931]  = 255;
  ram[7932]  = 255;
  ram[7933]  = 255;
  ram[7934]  = 255;
  ram[7935]  = 255;
  ram[7936]  = 255;
  ram[7937]  = 255;
  ram[7938]  = 255;
  ram[7939]  = 255;
  ram[7940]  = 255;
  ram[7941]  = 255;
  ram[7942]  = 255;
  ram[7943]  = 255;
  ram[7944]  = 255;
  ram[7945]  = 255;
  ram[7946]  = 255;
  ram[7947]  = 255;
  ram[7948]  = 255;
  ram[7949]  = 255;
  ram[7950]  = 255;
  ram[7951]  = 255;
  ram[7952]  = 255;
  ram[7953]  = 255;
  ram[7954]  = 255;
  ram[7955]  = 255;
  ram[7956]  = 255;
  ram[7957]  = 255;
  ram[7958]  = 255;
  ram[7959]  = 255;
  ram[7960]  = 255;
  ram[7961]  = 255;
  ram[7962]  = 255;
  ram[7963]  = 255;
  ram[7964]  = 255;
  ram[7965]  = 255;
  ram[7966]  = 255;
  ram[7967]  = 255;
  ram[7968]  = 255;
  ram[7969]  = 255;
  ram[7970]  = 255;
  ram[7971]  = 255;
  ram[7972]  = 255;
  ram[7973]  = 255;
  ram[7974]  = 255;
  ram[7975]  = 255;
  ram[7976]  = 255;
  ram[7977]  = 255;
  ram[7978]  = 255;
  ram[7979]  = 255;
  ram[7980]  = 255;
  ram[7981]  = 255;
  ram[7982]  = 255;
  ram[7983]  = 255;
  ram[7984]  = 255;
  ram[7985]  = 255;
  ram[7986]  = 255;
  ram[7987]  = 255;
  ram[7988]  = 255;
  ram[7989]  = 255;
  ram[7990]  = 255;
  ram[7991]  = 255;
  ram[7992]  = 255;
  ram[7993]  = 255;
  ram[7994]  = 255;
  ram[7995]  = 255;
  ram[7996]  = 236;
  ram[7997]  = 211;
  ram[7998]  = 243;
  ram[7999]  = 255;
  ram[8000]  = 255;
  ram[8001]  = 233;
  ram[8002]  = 204;
  ram[8003]  = 243;
  ram[8004]  = 255;
  ram[8005]  = 254;
  ram[8006]  = 251;
  ram[8007]  = 255;
  ram[8008]  = 255;
  ram[8009]  = 255;
  ram[8010]  = 255;
  ram[8011]  = 255;
  ram[8012]  = 255;
  ram[8013]  = 255;
  ram[8014]  = 255;
  ram[8015]  = 255;
  ram[8016]  = 255;
  ram[8017]  = 255;
  ram[8018]  = 255;
  ram[8019]  = 255;
  ram[8020]  = 255;
  ram[8021]  = 255;
  ram[8022]  = 255;
  ram[8023]  = 255;
  ram[8024]  = 255;
  ram[8025]  = 255;
  ram[8026]  = 255;
  ram[8027]  = 255;
  ram[8028]  = 255;
  ram[8029]  = 255;
  ram[8030]  = 255;
  ram[8031]  = 255;
  ram[8032]  = 255;
  ram[8033]  = 255;
  ram[8034]  = 255;
  ram[8035]  = 255;
  ram[8036]  = 255;
  ram[8037]  = 255;
  ram[8038]  = 255;
  ram[8039]  = 255;
  ram[8040]  = 255;
  ram[8041]  = 255;
  ram[8042]  = 255;
  ram[8043]  = 255;
  ram[8044]  = 255;
  ram[8045]  = 255;
  ram[8046]  = 255;
  ram[8047]  = 255;
  ram[8048]  = 255;
  ram[8049]  = 255;
  ram[8050]  = 255;
  ram[8051]  = 255;
  ram[8052]  = 255;
  ram[8053]  = 255;
  ram[8054]  = 255;
  ram[8055]  = 255;
  ram[8056]  = 255;
  ram[8057]  = 255;
  ram[8058]  = 255;
  ram[8059]  = 255;
  ram[8060]  = 255;
  ram[8061]  = 255;
  ram[8062]  = 255;
  ram[8063]  = 255;
  ram[8064]  = 255;
  ram[8065]  = 255;
  ram[8066]  = 255;
  ram[8067]  = 255;
  ram[8068]  = 255;
  ram[8069]  = 255;
  ram[8070]  = 255;
  ram[8071]  = 255;
  ram[8072]  = 255;
  ram[8073]  = 255;
  ram[8074]  = 255;
  ram[8075]  = 255;
  ram[8076]  = 255;
  ram[8077]  = 255;
  ram[8078]  = 255;
  ram[8079]  = 255;
  ram[8080]  = 255;
  ram[8081]  = 255;
  ram[8082]  = 255;
  ram[8083]  = 255;
  ram[8084]  = 255;
  ram[8085]  = 255;
  ram[8086]  = 255;
  ram[8087]  = 255;
  ram[8088]  = 255;
  ram[8089]  = 255;
  ram[8090]  = 255;
  ram[8091]  = 255;
  ram[8092]  = 255;
  ram[8093]  = 255;
  ram[8094]  = 255;
  ram[8095]  = 255;
  ram[8096]  = 255;
  ram[8097]  = 255;
  ram[8098]  = 255;
  ram[8099]  = 255;
  ram[8100]  = 255;
  ram[8101]  = 255;
  ram[8102]  = 255;
  ram[8103]  = 255;
  ram[8104]  = 255;
  ram[8105]  = 255;
  ram[8106]  = 255;
  ram[8107]  = 255;
  ram[8108]  = 255;
  ram[8109]  = 255;
  ram[8110]  = 255;
  ram[8111]  = 255;
  ram[8112]  = 255;
  ram[8113]  = 255;
  ram[8114]  = 255;
  ram[8115]  = 255;
  ram[8116]  = 255;
  ram[8117]  = 255;
  ram[8118]  = 255;
  ram[8119]  = 255;
  ram[8120]  = 255;
  ram[8121]  = 255;
  ram[8122]  = 255;
  ram[8123]  = 255;
  ram[8124]  = 255;
  ram[8125]  = 255;
  ram[8126]  = 255;
  ram[8127]  = 255;
  ram[8128]  = 255;
  ram[8129]  = 255;
  ram[8130]  = 255;
  ram[8131]  = 255;
  ram[8132]  = 255;
  ram[8133]  = 255;
  ram[8134]  = 255;
  ram[8135]  = 255;
  ram[8136]  = 255;
  ram[8137]  = 255;
  ram[8138]  = 255;
  ram[8139]  = 255;
  ram[8140]  = 255;
  ram[8141]  = 255;
  ram[8142]  = 255;
  ram[8143]  = 255;
  ram[8144]  = 255;
  ram[8145]  = 255;
  ram[8146]  = 255;
  ram[8147]  = 255;
  ram[8148]  = 255;
  ram[8149]  = 255;
  ram[8150]  = 255;
  ram[8151]  = 255;
  ram[8152]  = 255;
  ram[8153]  = 255;
  ram[8154]  = 255;
  ram[8155]  = 255;
  ram[8156]  = 255;
  ram[8157]  = 255;
  ram[8158]  = 255;
  ram[8159]  = 255;
  ram[8160]  = 255;
  ram[8161]  = 255;
  ram[8162]  = 255;
  ram[8163]  = 255;
  ram[8164]  = 255;
  ram[8165]  = 255;
  ram[8166]  = 255;
  ram[8167]  = 255;
  ram[8168]  = 255;
  ram[8169]  = 255;
  ram[8170]  = 255;
  ram[8171]  = 255;
  ram[8172]  = 255;
  ram[8173]  = 255;
  ram[8174]  = 255;
  ram[8175]  = 255;
  ram[8176]  = 255;
  ram[8177]  = 255;
  ram[8178]  = 255;
  ram[8179]  = 255;
  ram[8180]  = 255;
  ram[8181]  = 255;
  ram[8182]  = 255;
  ram[8183]  = 255;
  ram[8184]  = 255;
  ram[8185]  = 255;
  ram[8186]  = 255;
  ram[8187]  = 255;
  ram[8188]  = 255;
  ram[8189]  = 255;
  ram[8190]  = 255;
  ram[8191]  = 255;
  ram[8192]  = 255;
  ram[8193]  = 255;
  ram[8194]  = 255;
  ram[8195]  = 255;
  ram[8196]  = 236;
  ram[8197]  = 211;
  ram[8198]  = 243;
  ram[8199]  = 255;
  ram[8200]  = 255;
  ram[8201]  = 234;
  ram[8202]  = 204;
  ram[8203]  = 243;
  ram[8204]  = 254;
  ram[8205]  = 254;
  ram[8206]  = 250;
  ram[8207]  = 255;
  ram[8208]  = 255;
  ram[8209]  = 255;
  ram[8210]  = 255;
  ram[8211]  = 255;
  ram[8212]  = 255;
  ram[8213]  = 255;
  ram[8214]  = 255;
  ram[8215]  = 255;
  ram[8216]  = 255;
  ram[8217]  = 255;
  ram[8218]  = 255;
  ram[8219]  = 255;
  ram[8220]  = 255;
  ram[8221]  = 255;
  ram[8222]  = 255;
  ram[8223]  = 255;
  ram[8224]  = 255;
  ram[8225]  = 255;
  ram[8226]  = 255;
  ram[8227]  = 255;
  ram[8228]  = 255;
  ram[8229]  = 255;
  ram[8230]  = 255;
  ram[8231]  = 255;
  ram[8232]  = 255;
  ram[8233]  = 255;
  ram[8234]  = 255;
  ram[8235]  = 255;
  ram[8236]  = 255;
  ram[8237]  = 255;
  ram[8238]  = 255;
  ram[8239]  = 255;
  ram[8240]  = 255;
  ram[8241]  = 255;
  ram[8242]  = 255;
  ram[8243]  = 255;
  ram[8244]  = 255;
  ram[8245]  = 255;
  ram[8246]  = 255;
  ram[8247]  = 255;
  ram[8248]  = 255;
  ram[8249]  = 255;
  ram[8250]  = 255;
  ram[8251]  = 255;
  ram[8252]  = 255;
  ram[8253]  = 255;
  ram[8254]  = 255;
  ram[8255]  = 255;
  ram[8256]  = 255;
  ram[8257]  = 255;
  ram[8258]  = 255;
  ram[8259]  = 255;
  ram[8260]  = 255;
  ram[8261]  = 255;
  ram[8262]  = 255;
  ram[8263]  = 255;
  ram[8264]  = 255;
  ram[8265]  = 255;
  ram[8266]  = 255;
  ram[8267]  = 255;
  ram[8268]  = 255;
  ram[8269]  = 255;
  ram[8270]  = 255;
  ram[8271]  = 255;
  ram[8272]  = 255;
  ram[8273]  = 255;
  ram[8274]  = 255;
  ram[8275]  = 255;
  ram[8276]  = 255;
  ram[8277]  = 255;
  ram[8278]  = 255;
  ram[8279]  = 255;
  ram[8280]  = 255;
  ram[8281]  = 255;
  ram[8282]  = 255;
  ram[8283]  = 255;
  ram[8284]  = 255;
  ram[8285]  = 255;
  ram[8286]  = 255;
  ram[8287]  = 255;
  ram[8288]  = 255;
  ram[8289]  = 255;
  ram[8290]  = 255;
  ram[8291]  = 255;
  ram[8292]  = 255;
  ram[8293]  = 255;
  ram[8294]  = 255;
  ram[8295]  = 255;
  ram[8296]  = 255;
  ram[8297]  = 255;
  ram[8298]  = 255;
  ram[8299]  = 255;
  ram[8300]  = 255;
  ram[8301]  = 255;
  ram[8302]  = 255;
  ram[8303]  = 255;
  ram[8304]  = 255;
  ram[8305]  = 255;
  ram[8306]  = 255;
  ram[8307]  = 255;
  ram[8308]  = 255;
  ram[8309]  = 255;
  ram[8310]  = 255;
  ram[8311]  = 255;
  ram[8312]  = 255;
  ram[8313]  = 255;
  ram[8314]  = 255;
  ram[8315]  = 255;
  ram[8316]  = 255;
  ram[8317]  = 255;
  ram[8318]  = 255;
  ram[8319]  = 255;
  ram[8320]  = 255;
  ram[8321]  = 255;
  ram[8322]  = 255;
  ram[8323]  = 255;
  ram[8324]  = 255;
  ram[8325]  = 255;
  ram[8326]  = 255;
  ram[8327]  = 255;
  ram[8328]  = 255;
  ram[8329]  = 255;
  ram[8330]  = 255;
  ram[8331]  = 255;
  ram[8332]  = 255;
  ram[8333]  = 255;
  ram[8334]  = 255;
  ram[8335]  = 255;
  ram[8336]  = 255;
  ram[8337]  = 255;
  ram[8338]  = 255;
  ram[8339]  = 255;
  ram[8340]  = 255;
  ram[8341]  = 255;
  ram[8342]  = 255;
  ram[8343]  = 255;
  ram[8344]  = 255;
  ram[8345]  = 255;
  ram[8346]  = 255;
  ram[8347]  = 255;
  ram[8348]  = 255;
  ram[8349]  = 255;
  ram[8350]  = 255;
  ram[8351]  = 255;
  ram[8352]  = 255;
  ram[8353]  = 255;
  ram[8354]  = 255;
  ram[8355]  = 255;
  ram[8356]  = 255;
  ram[8357]  = 255;
  ram[8358]  = 255;
  ram[8359]  = 255;
  ram[8360]  = 255;
  ram[8361]  = 255;
  ram[8362]  = 255;
  ram[8363]  = 255;
  ram[8364]  = 255;
  ram[8365]  = 255;
  ram[8366]  = 255;
  ram[8367]  = 255;
  ram[8368]  = 255;
  ram[8369]  = 255;
  ram[8370]  = 255;
  ram[8371]  = 255;
  ram[8372]  = 255;
  ram[8373]  = 255;
  ram[8374]  = 255;
  ram[8375]  = 255;
  ram[8376]  = 255;
  ram[8377]  = 255;
  ram[8378]  = 255;
  ram[8379]  = 255;
  ram[8380]  = 255;
  ram[8381]  = 255;
  ram[8382]  = 255;
  ram[8383]  = 255;
  ram[8384]  = 255;
  ram[8385]  = 255;
  ram[8386]  = 255;
  ram[8387]  = 255;
  ram[8388]  = 255;
  ram[8389]  = 255;
  ram[8390]  = 255;
  ram[8391]  = 255;
  ram[8392]  = 255;
  ram[8393]  = 255;
  ram[8394]  = 255;
  ram[8395]  = 255;
  ram[8396]  = 236;
  ram[8397]  = 211;
  ram[8398]  = 243;
  ram[8399]  = 255;
  ram[8400]  = 255;
  ram[8401]  = 234;
  ram[8402]  = 205;
  ram[8403]  = 243;
  ram[8404]  = 255;
  ram[8405]  = 254;
  ram[8406]  = 250;
  ram[8407]  = 255;
  ram[8408]  = 255;
  ram[8409]  = 255;
  ram[8410]  = 255;
  ram[8411]  = 255;
  ram[8412]  = 255;
  ram[8413]  = 255;
  ram[8414]  = 255;
  ram[8415]  = 255;
  ram[8416]  = 255;
  ram[8417]  = 255;
  ram[8418]  = 255;
  ram[8419]  = 255;
  ram[8420]  = 255;
  ram[8421]  = 255;
  ram[8422]  = 255;
  ram[8423]  = 255;
  ram[8424]  = 255;
  ram[8425]  = 255;
  ram[8426]  = 255;
  ram[8427]  = 255;
  ram[8428]  = 255;
  ram[8429]  = 255;
  ram[8430]  = 255;
  ram[8431]  = 255;
  ram[8432]  = 255;
  ram[8433]  = 255;
  ram[8434]  = 255;
  ram[8435]  = 255;
  ram[8436]  = 255;
  ram[8437]  = 255;
  ram[8438]  = 255;
  ram[8439]  = 255;
  ram[8440]  = 255;
  ram[8441]  = 255;
  ram[8442]  = 255;
  ram[8443]  = 255;
  ram[8444]  = 255;
  ram[8445]  = 255;
  ram[8446]  = 255;
  ram[8447]  = 255;
  ram[8448]  = 255;
  ram[8449]  = 255;
  ram[8450]  = 255;
  ram[8451]  = 255;
  ram[8452]  = 255;
  ram[8453]  = 255;
  ram[8454]  = 255;
  ram[8455]  = 255;
  ram[8456]  = 255;
  ram[8457]  = 255;
  ram[8458]  = 255;
  ram[8459]  = 255;
  ram[8460]  = 255;
  ram[8461]  = 255;
  ram[8462]  = 255;
  ram[8463]  = 255;
  ram[8464]  = 255;
  ram[8465]  = 255;
  ram[8466]  = 255;
  ram[8467]  = 255;
  ram[8468]  = 255;
  ram[8469]  = 255;
  ram[8470]  = 255;
  ram[8471]  = 255;
  ram[8472]  = 255;
  ram[8473]  = 255;
  ram[8474]  = 255;
  ram[8475]  = 255;
  ram[8476]  = 255;
  ram[8477]  = 255;
  ram[8478]  = 255;
  ram[8479]  = 255;
  ram[8480]  = 255;
  ram[8481]  = 255;
  ram[8482]  = 255;
  ram[8483]  = 255;
  ram[8484]  = 255;
  ram[8485]  = 255;
  ram[8486]  = 255;
  ram[8487]  = 255;
  ram[8488]  = 255;
  ram[8489]  = 255;
  ram[8490]  = 255;
  ram[8491]  = 255;
  ram[8492]  = 255;
  ram[8493]  = 255;
  ram[8494]  = 255;
  ram[8495]  = 255;
  ram[8496]  = 255;
  ram[8497]  = 255;
  ram[8498]  = 255;
  ram[8499]  = 255;
  ram[8500]  = 255;
  ram[8501]  = 255;
  ram[8502]  = 255;
  ram[8503]  = 255;
  ram[8504]  = 255;
  ram[8505]  = 255;
  ram[8506]  = 255;
  ram[8507]  = 255;
  ram[8508]  = 255;
  ram[8509]  = 255;
  ram[8510]  = 255;
  ram[8511]  = 255;
  ram[8512]  = 255;
  ram[8513]  = 255;
  ram[8514]  = 255;
  ram[8515]  = 255;
  ram[8516]  = 255;
  ram[8517]  = 255;
  ram[8518]  = 255;
  ram[8519]  = 255;
  ram[8520]  = 255;
  ram[8521]  = 255;
  ram[8522]  = 255;
  ram[8523]  = 255;
  ram[8524]  = 255;
  ram[8525]  = 255;
  ram[8526]  = 255;
  ram[8527]  = 255;
  ram[8528]  = 255;
  ram[8529]  = 255;
  ram[8530]  = 255;
  ram[8531]  = 255;
  ram[8532]  = 255;
  ram[8533]  = 255;
  ram[8534]  = 255;
  ram[8535]  = 255;
  ram[8536]  = 255;
  ram[8537]  = 255;
  ram[8538]  = 255;
  ram[8539]  = 255;
  ram[8540]  = 255;
  ram[8541]  = 255;
  ram[8542]  = 255;
  ram[8543]  = 255;
  ram[8544]  = 255;
  ram[8545]  = 255;
  ram[8546]  = 255;
  ram[8547]  = 255;
  ram[8548]  = 255;
  ram[8549]  = 255;
  ram[8550]  = 255;
  ram[8551]  = 255;
  ram[8552]  = 255;
  ram[8553]  = 255;
  ram[8554]  = 255;
  ram[8555]  = 255;
  ram[8556]  = 255;
  ram[8557]  = 255;
  ram[8558]  = 255;
  ram[8559]  = 255;
  ram[8560]  = 255;
  ram[8561]  = 255;
  ram[8562]  = 255;
  ram[8563]  = 255;
  ram[8564]  = 255;
  ram[8565]  = 255;
  ram[8566]  = 255;
  ram[8567]  = 255;
  ram[8568]  = 255;
  ram[8569]  = 255;
  ram[8570]  = 255;
  ram[8571]  = 255;
  ram[8572]  = 255;
  ram[8573]  = 255;
  ram[8574]  = 255;
  ram[8575]  = 255;
  ram[8576]  = 255;
  ram[8577]  = 255;
  ram[8578]  = 255;
  ram[8579]  = 255;
  ram[8580]  = 255;
  ram[8581]  = 255;
  ram[8582]  = 255;
  ram[8583]  = 255;
  ram[8584]  = 255;
  ram[8585]  = 255;
  ram[8586]  = 255;
  ram[8587]  = 255;
  ram[8588]  = 255;
  ram[8589]  = 255;
  ram[8590]  = 255;
  ram[8591]  = 255;
  ram[8592]  = 255;
  ram[8593]  = 255;
  ram[8594]  = 255;
  ram[8595]  = 255;
  ram[8596]  = 236;
  ram[8597]  = 211;
  ram[8598]  = 243;
  ram[8599]  = 255;
  ram[8600]  = 255;
  ram[8601]  = 234;
  ram[8602]  = 206;
  ram[8603]  = 243;
  ram[8604]  = 255;
  ram[8605]  = 254;
  ram[8606]  = 251;
  ram[8607]  = 255;
  ram[8608]  = 255;
  ram[8609]  = 255;
  ram[8610]  = 255;
  ram[8611]  = 255;
  ram[8612]  = 255;
  ram[8613]  = 255;
  ram[8614]  = 255;
  ram[8615]  = 255;
  ram[8616]  = 255;
  ram[8617]  = 255;
  ram[8618]  = 255;
  ram[8619]  = 255;
  ram[8620]  = 255;
  ram[8621]  = 255;
  ram[8622]  = 255;
  ram[8623]  = 255;
  ram[8624]  = 255;
  ram[8625]  = 255;
  ram[8626]  = 255;
  ram[8627]  = 255;
  ram[8628]  = 255;
  ram[8629]  = 255;
  ram[8630]  = 255;
  ram[8631]  = 255;
  ram[8632]  = 255;
  ram[8633]  = 255;
  ram[8634]  = 255;
  ram[8635]  = 255;
  ram[8636]  = 255;
  ram[8637]  = 255;
  ram[8638]  = 255;
  ram[8639]  = 255;
  ram[8640]  = 255;
  ram[8641]  = 255;
  ram[8642]  = 255;
  ram[8643]  = 255;
  ram[8644]  = 255;
  ram[8645]  = 255;
  ram[8646]  = 255;
  ram[8647]  = 255;
  ram[8648]  = 255;
  ram[8649]  = 255;
  ram[8650]  = 255;
  ram[8651]  = 255;
  ram[8652]  = 255;
  ram[8653]  = 255;
  ram[8654]  = 255;
  ram[8655]  = 255;
  ram[8656]  = 255;
  ram[8657]  = 255;
  ram[8658]  = 255;
  ram[8659]  = 255;
  ram[8660]  = 255;
  ram[8661]  = 255;
  ram[8662]  = 255;
  ram[8663]  = 255;
  ram[8664]  = 255;
  ram[8665]  = 255;
  ram[8666]  = 255;
  ram[8667]  = 255;
  ram[8668]  = 255;
  ram[8669]  = 255;
  ram[8670]  = 255;
  ram[8671]  = 255;
  ram[8672]  = 255;
  ram[8673]  = 255;
  ram[8674]  = 255;
  ram[8675]  = 255;
  ram[8676]  = 255;
  ram[8677]  = 255;
  ram[8678]  = 255;
  ram[8679]  = 255;
  ram[8680]  = 255;
  ram[8681]  = 255;
  ram[8682]  = 255;
  ram[8683]  = 255;
  ram[8684]  = 255;
  ram[8685]  = 255;
  ram[8686]  = 255;
  ram[8687]  = 255;
  ram[8688]  = 255;
  ram[8689]  = 255;
  ram[8690]  = 255;
  ram[8691]  = 255;
  ram[8692]  = 255;
  ram[8693]  = 255;
  ram[8694]  = 255;
  ram[8695]  = 255;
  ram[8696]  = 255;
  ram[8697]  = 255;
  ram[8698]  = 255;
  ram[8699]  = 255;
  ram[8700]  = 255;
  ram[8701]  = 255;
  ram[8702]  = 255;
  ram[8703]  = 255;
  ram[8704]  = 255;
  ram[8705]  = 255;
  ram[8706]  = 255;
  ram[8707]  = 255;
  ram[8708]  = 255;
  ram[8709]  = 255;
  ram[8710]  = 255;
  ram[8711]  = 255;
  ram[8712]  = 255;
  ram[8713]  = 255;
  ram[8714]  = 255;
  ram[8715]  = 255;
  ram[8716]  = 255;
  ram[8717]  = 255;
  ram[8718]  = 255;
  ram[8719]  = 255;
  ram[8720]  = 255;
  ram[8721]  = 255;
  ram[8722]  = 255;
  ram[8723]  = 255;
  ram[8724]  = 255;
  ram[8725]  = 255;
  ram[8726]  = 255;
  ram[8727]  = 255;
  ram[8728]  = 255;
  ram[8729]  = 255;
  ram[8730]  = 255;
  ram[8731]  = 255;
  ram[8732]  = 255;
  ram[8733]  = 255;
  ram[8734]  = 255;
  ram[8735]  = 255;
  ram[8736]  = 255;
  ram[8737]  = 255;
  ram[8738]  = 255;
  ram[8739]  = 255;
  ram[8740]  = 255;
  ram[8741]  = 255;
  ram[8742]  = 255;
  ram[8743]  = 255;
  ram[8744]  = 255;
  ram[8745]  = 255;
  ram[8746]  = 255;
  ram[8747]  = 255;
  ram[8748]  = 255;
  ram[8749]  = 255;
  ram[8750]  = 255;
  ram[8751]  = 255;
  ram[8752]  = 255;
  ram[8753]  = 255;
  ram[8754]  = 255;
  ram[8755]  = 255;
  ram[8756]  = 255;
  ram[8757]  = 255;
  ram[8758]  = 255;
  ram[8759]  = 255;
  ram[8760]  = 255;
  ram[8761]  = 255;
  ram[8762]  = 255;
  ram[8763]  = 255;
  ram[8764]  = 255;
  ram[8765]  = 255;
  ram[8766]  = 255;
  ram[8767]  = 255;
  ram[8768]  = 255;
  ram[8769]  = 255;
  ram[8770]  = 255;
  ram[8771]  = 255;
  ram[8772]  = 255;
  ram[8773]  = 255;
  ram[8774]  = 255;
  ram[8775]  = 255;
  ram[8776]  = 255;
  ram[8777]  = 255;
  ram[8778]  = 255;
  ram[8779]  = 255;
  ram[8780]  = 255;
  ram[8781]  = 255;
  ram[8782]  = 255;
  ram[8783]  = 255;
  ram[8784]  = 255;
  ram[8785]  = 255;
  ram[8786]  = 255;
  ram[8787]  = 255;
  ram[8788]  = 255;
  ram[8789]  = 255;
  ram[8790]  = 255;
  ram[8791]  = 255;
  ram[8792]  = 255;
  ram[8793]  = 255;
  ram[8794]  = 255;
  ram[8795]  = 255;
  ram[8796]  = 236;
  ram[8797]  = 212;
  ram[8798]  = 243;
  ram[8799]  = 255;
  ram[8800]  = 255;
  ram[8801]  = 233;
  ram[8802]  = 194;
  ram[8803]  = 242;
  ram[8804]  = 255;
  ram[8805]  = 255;
  ram[8806]  = 255;
  ram[8807]  = 255;
  ram[8808]  = 255;
  ram[8809]  = 255;
  ram[8810]  = 255;
  ram[8811]  = 255;
  ram[8812]  = 255;
  ram[8813]  = 255;
  ram[8814]  = 255;
  ram[8815]  = 255;
  ram[8816]  = 255;
  ram[8817]  = 255;
  ram[8818]  = 255;
  ram[8819]  = 255;
  ram[8820]  = 255;
  ram[8821]  = 255;
  ram[8822]  = 255;
  ram[8823]  = 255;
  ram[8824]  = 255;
  ram[8825]  = 255;
  ram[8826]  = 255;
  ram[8827]  = 255;
  ram[8828]  = 255;
  ram[8829]  = 255;
  ram[8830]  = 255;
  ram[8831]  = 255;
  ram[8832]  = 255;
  ram[8833]  = 255;
  ram[8834]  = 255;
  ram[8835]  = 255;
  ram[8836]  = 255;
  ram[8837]  = 255;
  ram[8838]  = 255;
  ram[8839]  = 255;
  ram[8840]  = 255;
  ram[8841]  = 255;
  ram[8842]  = 255;
  ram[8843]  = 255;
  ram[8844]  = 255;
  ram[8845]  = 255;
  ram[8846]  = 255;
  ram[8847]  = 255;
  ram[8848]  = 255;
  ram[8849]  = 255;
  ram[8850]  = 255;
  ram[8851]  = 255;
  ram[8852]  = 255;
  ram[8853]  = 255;
  ram[8854]  = 255;
  ram[8855]  = 255;
  ram[8856]  = 255;
  ram[8857]  = 255;
  ram[8858]  = 255;
  ram[8859]  = 255;
  ram[8860]  = 255;
  ram[8861]  = 255;
  ram[8862]  = 255;
  ram[8863]  = 255;
  ram[8864]  = 255;
  ram[8865]  = 255;
  ram[8866]  = 255;
  ram[8867]  = 255;
  ram[8868]  = 255;
  ram[8869]  = 255;
  ram[8870]  = 255;
  ram[8871]  = 255;
  ram[8872]  = 255;
  ram[8873]  = 255;
  ram[8874]  = 255;
  ram[8875]  = 255;
  ram[8876]  = 255;
  ram[8877]  = 255;
  ram[8878]  = 255;
  ram[8879]  = 255;
  ram[8880]  = 255;
  ram[8881]  = 255;
  ram[8882]  = 255;
  ram[8883]  = 255;
  ram[8884]  = 255;
  ram[8885]  = 255;
  ram[8886]  = 255;
  ram[8887]  = 255;
  ram[8888]  = 255;
  ram[8889]  = 255;
  ram[8890]  = 255;
  ram[8891]  = 255;
  ram[8892]  = 255;
  ram[8893]  = 255;
  ram[8894]  = 255;
  ram[8895]  = 255;
  ram[8896]  = 255;
  ram[8897]  = 255;
  ram[8898]  = 255;
  ram[8899]  = 255;
  ram[8900]  = 255;
  ram[8901]  = 255;
  ram[8902]  = 255;
  ram[8903]  = 255;
  ram[8904]  = 255;
  ram[8905]  = 255;
  ram[8906]  = 255;
  ram[8907]  = 255;
  ram[8908]  = 255;
  ram[8909]  = 255;
  ram[8910]  = 255;
  ram[8911]  = 255;
  ram[8912]  = 255;
  ram[8913]  = 255;
  ram[8914]  = 255;
  ram[8915]  = 255;
  ram[8916]  = 255;
  ram[8917]  = 255;
  ram[8918]  = 255;
  ram[8919]  = 255;
  ram[8920]  = 255;
  ram[8921]  = 255;
  ram[8922]  = 255;
  ram[8923]  = 255;
  ram[8924]  = 255;
  ram[8925]  = 255;
  ram[8926]  = 255;
  ram[8927]  = 255;
  ram[8928]  = 255;
  ram[8929]  = 255;
  ram[8930]  = 255;
  ram[8931]  = 255;
  ram[8932]  = 255;
  ram[8933]  = 255;
  ram[8934]  = 255;
  ram[8935]  = 255;
  ram[8936]  = 255;
  ram[8937]  = 255;
  ram[8938]  = 255;
  ram[8939]  = 255;
  ram[8940]  = 255;
  ram[8941]  = 255;
  ram[8942]  = 255;
  ram[8943]  = 255;
  ram[8944]  = 255;
  ram[8945]  = 255;
  ram[8946]  = 255;
  ram[8947]  = 255;
  ram[8948]  = 255;
  ram[8949]  = 255;
  ram[8950]  = 255;
  ram[8951]  = 255;
  ram[8952]  = 255;
  ram[8953]  = 255;
  ram[8954]  = 255;
  ram[8955]  = 255;
  ram[8956]  = 255;
  ram[8957]  = 255;
  ram[8958]  = 255;
  ram[8959]  = 255;
  ram[8960]  = 255;
  ram[8961]  = 255;
  ram[8962]  = 255;
  ram[8963]  = 255;
  ram[8964]  = 255;
  ram[8965]  = 255;
  ram[8966]  = 255;
  ram[8967]  = 255;
  ram[8968]  = 255;
  ram[8969]  = 255;
  ram[8970]  = 255;
  ram[8971]  = 255;
  ram[8972]  = 255;
  ram[8973]  = 255;
  ram[8974]  = 255;
  ram[8975]  = 255;
  ram[8976]  = 255;
  ram[8977]  = 255;
  ram[8978]  = 255;
  ram[8979]  = 255;
  ram[8980]  = 255;
  ram[8981]  = 255;
  ram[8982]  = 255;
  ram[8983]  = 255;
  ram[8984]  = 255;
  ram[8985]  = 255;
  ram[8986]  = 255;
  ram[8987]  = 255;
  ram[8988]  = 255;
  ram[8989]  = 255;
  ram[8990]  = 255;
  ram[8991]  = 255;
  ram[8992]  = 255;
  ram[8993]  = 255;
  ram[8994]  = 255;
  ram[8995]  = 255;
  ram[8996]  = 233;
  ram[8997]  = 202;
  ram[8998]  = 239;
  ram[8999]  = 255;
  ram[9000]  = 255;
  ram[9001]  = 233;
  ram[9002]  = 211;
  ram[9003]  = 236;
  ram[9004]  = 225;
  ram[9005]  = 223;
  ram[9006]  = 228;
  ram[9007]  = 229;
  ram[9008]  = 229;
  ram[9009]  = 229;
  ram[9010]  = 229;
  ram[9011]  = 229;
  ram[9012]  = 229;
  ram[9013]  = 229;
  ram[9014]  = 229;
  ram[9015]  = 229;
  ram[9016]  = 229;
  ram[9017]  = 229;
  ram[9018]  = 229;
  ram[9019]  = 229;
  ram[9020]  = 229;
  ram[9021]  = 229;
  ram[9022]  = 229;
  ram[9023]  = 229;
  ram[9024]  = 230;
  ram[9025]  = 230;
  ram[9026]  = 230;
  ram[9027]  = 230;
  ram[9028]  = 230;
  ram[9029]  = 230;
  ram[9030]  = 230;
  ram[9031]  = 230;
  ram[9032]  = 230;
  ram[9033]  = 230;
  ram[9034]  = 230;
  ram[9035]  = 230;
  ram[9036]  = 230;
  ram[9037]  = 230;
  ram[9038]  = 230;
  ram[9039]  = 230;
  ram[9040]  = 230;
  ram[9041]  = 230;
  ram[9042]  = 230;
  ram[9043]  = 230;
  ram[9044]  = 230;
  ram[9045]  = 230;
  ram[9046]  = 230;
  ram[9047]  = 230;
  ram[9048]  = 230;
  ram[9049]  = 230;
  ram[9050]  = 230;
  ram[9051]  = 230;
  ram[9052]  = 230;
  ram[9053]  = 230;
  ram[9054]  = 230;
  ram[9055]  = 230;
  ram[9056]  = 230;
  ram[9057]  = 230;
  ram[9058]  = 230;
  ram[9059]  = 230;
  ram[9060]  = 230;
  ram[9061]  = 230;
  ram[9062]  = 230;
  ram[9063]  = 230;
  ram[9064]  = 230;
  ram[9065]  = 230;
  ram[9066]  = 230;
  ram[9067]  = 230;
  ram[9068]  = 230;
  ram[9069]  = 230;
  ram[9070]  = 230;
  ram[9071]  = 230;
  ram[9072]  = 230;
  ram[9073]  = 230;
  ram[9074]  = 230;
  ram[9075]  = 230;
  ram[9076]  = 230;
  ram[9077]  = 230;
  ram[9078]  = 230;
  ram[9079]  = 230;
  ram[9080]  = 230;
  ram[9081]  = 230;
  ram[9082]  = 230;
  ram[9083]  = 230;
  ram[9084]  = 230;
  ram[9085]  = 230;
  ram[9086]  = 230;
  ram[9087]  = 230;
  ram[9088]  = 230;
  ram[9089]  = 230;
  ram[9090]  = 230;
  ram[9091]  = 230;
  ram[9092]  = 230;
  ram[9093]  = 230;
  ram[9094]  = 230;
  ram[9095]  = 230;
  ram[9096]  = 230;
  ram[9097]  = 230;
  ram[9098]  = 230;
  ram[9099]  = 230;
  ram[9100]  = 230;
  ram[9101]  = 230;
  ram[9102]  = 230;
  ram[9103]  = 230;
  ram[9104]  = 230;
  ram[9105]  = 230;
  ram[9106]  = 230;
  ram[9107]  = 230;
  ram[9108]  = 230;
  ram[9109]  = 230;
  ram[9110]  = 230;
  ram[9111]  = 230;
  ram[9112]  = 230;
  ram[9113]  = 230;
  ram[9114]  = 230;
  ram[9115]  = 230;
  ram[9116]  = 230;
  ram[9117]  = 230;
  ram[9118]  = 230;
  ram[9119]  = 230;
  ram[9120]  = 230;
  ram[9121]  = 230;
  ram[9122]  = 230;
  ram[9123]  = 230;
  ram[9124]  = 230;
  ram[9125]  = 230;
  ram[9126]  = 230;
  ram[9127]  = 230;
  ram[9128]  = 230;
  ram[9129]  = 230;
  ram[9130]  = 230;
  ram[9131]  = 230;
  ram[9132]  = 230;
  ram[9133]  = 230;
  ram[9134]  = 230;
  ram[9135]  = 230;
  ram[9136]  = 230;
  ram[9137]  = 230;
  ram[9138]  = 230;
  ram[9139]  = 230;
  ram[9140]  = 230;
  ram[9141]  = 230;
  ram[9142]  = 230;
  ram[9143]  = 230;
  ram[9144]  = 230;
  ram[9145]  = 230;
  ram[9146]  = 230;
  ram[9147]  = 230;
  ram[9148]  = 230;
  ram[9149]  = 230;
  ram[9150]  = 230;
  ram[9151]  = 230;
  ram[9152]  = 230;
  ram[9153]  = 230;
  ram[9154]  = 230;
  ram[9155]  = 230;
  ram[9156]  = 230;
  ram[9157]  = 230;
  ram[9158]  = 230;
  ram[9159]  = 230;
  ram[9160]  = 230;
  ram[9161]  = 230;
  ram[9162]  = 230;
  ram[9163]  = 230;
  ram[9164]  = 230;
  ram[9165]  = 230;
  ram[9166]  = 230;
  ram[9167]  = 230;
  ram[9168]  = 230;
  ram[9169]  = 230;
  ram[9170]  = 230;
  ram[9171]  = 230;
  ram[9172]  = 230;
  ram[9173]  = 230;
  ram[9174]  = 230;
  ram[9175]  = 230;
  ram[9176]  = 230;
  ram[9177]  = 230;
  ram[9178]  = 230;
  ram[9179]  = 230;
  ram[9180]  = 230;
  ram[9181]  = 230;
  ram[9182]  = 230;
  ram[9183]  = 230;
  ram[9184]  = 230;
  ram[9185]  = 230;
  ram[9186]  = 230;
  ram[9187]  = 230;
  ram[9188]  = 230;
  ram[9189]  = 230;
  ram[9190]  = 230;
  ram[9191]  = 230;
  ram[9192]  = 230;
  ram[9193]  = 230;
  ram[9194]  = 231;
  ram[9195]  = 230;
  ram[9196]  = 229;
  ram[9197]  = 210;
  ram[9198]  = 240;
  ram[9199]  = 255;
  ram[9200]  = 255;
  ram[9201]  = 230;
  ram[9202]  = 219;
  ram[9203]  = 224;
  ram[9204]  = 213;
  ram[9205]  = 216;
  ram[9206]  = 224;
  ram[9207]  = 229;
  ram[9208]  = 228;
  ram[9209]  = 228;
  ram[9210]  = 228;
  ram[9211]  = 228;
  ram[9212]  = 228;
  ram[9213]  = 228;
  ram[9214]  = 228;
  ram[9215]  = 228;
  ram[9216]  = 228;
  ram[9217]  = 228;
  ram[9218]  = 228;
  ram[9219]  = 228;
  ram[9220]  = 228;
  ram[9221]  = 228;
  ram[9222]  = 229;
  ram[9223]  = 229;
  ram[9224]  = 228;
  ram[9225]  = 227;
  ram[9226]  = 227;
  ram[9227]  = 227;
  ram[9228]  = 227;
  ram[9229]  = 227;
  ram[9230]  = 227;
  ram[9231]  = 227;
  ram[9232]  = 227;
  ram[9233]  = 227;
  ram[9234]  = 227;
  ram[9235]  = 227;
  ram[9236]  = 227;
  ram[9237]  = 227;
  ram[9238]  = 227;
  ram[9239]  = 227;
  ram[9240]  = 227;
  ram[9241]  = 227;
  ram[9242]  = 227;
  ram[9243]  = 227;
  ram[9244]  = 227;
  ram[9245]  = 227;
  ram[9246]  = 227;
  ram[9247]  = 227;
  ram[9248]  = 227;
  ram[9249]  = 227;
  ram[9250]  = 227;
  ram[9251]  = 227;
  ram[9252]  = 227;
  ram[9253]  = 227;
  ram[9254]  = 227;
  ram[9255]  = 227;
  ram[9256]  = 227;
  ram[9257]  = 227;
  ram[9258]  = 227;
  ram[9259]  = 227;
  ram[9260]  = 227;
  ram[9261]  = 227;
  ram[9262]  = 227;
  ram[9263]  = 227;
  ram[9264]  = 227;
  ram[9265]  = 227;
  ram[9266]  = 227;
  ram[9267]  = 227;
  ram[9268]  = 227;
  ram[9269]  = 227;
  ram[9270]  = 227;
  ram[9271]  = 227;
  ram[9272]  = 227;
  ram[9273]  = 227;
  ram[9274]  = 227;
  ram[9275]  = 227;
  ram[9276]  = 227;
  ram[9277]  = 227;
  ram[9278]  = 227;
  ram[9279]  = 227;
  ram[9280]  = 227;
  ram[9281]  = 227;
  ram[9282]  = 227;
  ram[9283]  = 227;
  ram[9284]  = 227;
  ram[9285]  = 227;
  ram[9286]  = 227;
  ram[9287]  = 227;
  ram[9288]  = 227;
  ram[9289]  = 227;
  ram[9290]  = 227;
  ram[9291]  = 227;
  ram[9292]  = 227;
  ram[9293]  = 227;
  ram[9294]  = 227;
  ram[9295]  = 227;
  ram[9296]  = 227;
  ram[9297]  = 227;
  ram[9298]  = 227;
  ram[9299]  = 227;
  ram[9300]  = 227;
  ram[9301]  = 227;
  ram[9302]  = 227;
  ram[9303]  = 227;
  ram[9304]  = 227;
  ram[9305]  = 227;
  ram[9306]  = 227;
  ram[9307]  = 227;
  ram[9308]  = 227;
  ram[9309]  = 227;
  ram[9310]  = 227;
  ram[9311]  = 227;
  ram[9312]  = 227;
  ram[9313]  = 227;
  ram[9314]  = 227;
  ram[9315]  = 227;
  ram[9316]  = 227;
  ram[9317]  = 227;
  ram[9318]  = 227;
  ram[9319]  = 227;
  ram[9320]  = 227;
  ram[9321]  = 227;
  ram[9322]  = 227;
  ram[9323]  = 227;
  ram[9324]  = 227;
  ram[9325]  = 227;
  ram[9326]  = 227;
  ram[9327]  = 227;
  ram[9328]  = 227;
  ram[9329]  = 227;
  ram[9330]  = 227;
  ram[9331]  = 227;
  ram[9332]  = 227;
  ram[9333]  = 227;
  ram[9334]  = 227;
  ram[9335]  = 227;
  ram[9336]  = 227;
  ram[9337]  = 227;
  ram[9338]  = 227;
  ram[9339]  = 227;
  ram[9340]  = 227;
  ram[9341]  = 227;
  ram[9342]  = 227;
  ram[9343]  = 227;
  ram[9344]  = 227;
  ram[9345]  = 227;
  ram[9346]  = 227;
  ram[9347]  = 227;
  ram[9348]  = 227;
  ram[9349]  = 227;
  ram[9350]  = 227;
  ram[9351]  = 227;
  ram[9352]  = 227;
  ram[9353]  = 227;
  ram[9354]  = 227;
  ram[9355]  = 227;
  ram[9356]  = 227;
  ram[9357]  = 227;
  ram[9358]  = 227;
  ram[9359]  = 227;
  ram[9360]  = 227;
  ram[9361]  = 227;
  ram[9362]  = 227;
  ram[9363]  = 227;
  ram[9364]  = 227;
  ram[9365]  = 227;
  ram[9366]  = 227;
  ram[9367]  = 227;
  ram[9368]  = 227;
  ram[9369]  = 227;
  ram[9370]  = 227;
  ram[9371]  = 227;
  ram[9372]  = 227;
  ram[9373]  = 227;
  ram[9374]  = 227;
  ram[9375]  = 227;
  ram[9376]  = 227;
  ram[9377]  = 227;
  ram[9378]  = 227;
  ram[9379]  = 227;
  ram[9380]  = 227;
  ram[9381]  = 227;
  ram[9382]  = 227;
  ram[9383]  = 227;
  ram[9384]  = 227;
  ram[9385]  = 227;
  ram[9386]  = 227;
  ram[9387]  = 227;
  ram[9388]  = 227;
  ram[9389]  = 227;
  ram[9390]  = 227;
  ram[9391]  = 227;
  ram[9392]  = 227;
  ram[9393]  = 226;
  ram[9394]  = 227;
  ram[9395]  = 221;
  ram[9396]  = 221;
  ram[9397]  = 225;
  ram[9398]  = 246;
  ram[9399]  = 255;
  ram[9400]  = 252;
  ram[9401]  = 240;
  ram[9402]  = 197;
  ram[9403]  = 207;
  ram[9404]  = 213;
  ram[9405]  = 214;
  ram[9406]  = 214;
  ram[9407]  = 210;
  ram[9408]  = 210;
  ram[9409]  = 210;
  ram[9410]  = 210;
  ram[9411]  = 210;
  ram[9412]  = 210;
  ram[9413]  = 210;
  ram[9414]  = 210;
  ram[9415]  = 210;
  ram[9416]  = 210;
  ram[9417]  = 210;
  ram[9418]  = 210;
  ram[9419]  = 210;
  ram[9420]  = 210;
  ram[9421]  = 210;
  ram[9422]  = 209;
  ram[9423]  = 209;
  ram[9424]  = 210;
  ram[9425]  = 211;
  ram[9426]  = 211;
  ram[9427]  = 211;
  ram[9428]  = 211;
  ram[9429]  = 211;
  ram[9430]  = 211;
  ram[9431]  = 211;
  ram[9432]  = 211;
  ram[9433]  = 211;
  ram[9434]  = 211;
  ram[9435]  = 211;
  ram[9436]  = 211;
  ram[9437]  = 211;
  ram[9438]  = 211;
  ram[9439]  = 211;
  ram[9440]  = 211;
  ram[9441]  = 211;
  ram[9442]  = 211;
  ram[9443]  = 211;
  ram[9444]  = 211;
  ram[9445]  = 211;
  ram[9446]  = 211;
  ram[9447]  = 211;
  ram[9448]  = 211;
  ram[9449]  = 211;
  ram[9450]  = 211;
  ram[9451]  = 211;
  ram[9452]  = 211;
  ram[9453]  = 211;
  ram[9454]  = 211;
  ram[9455]  = 211;
  ram[9456]  = 211;
  ram[9457]  = 211;
  ram[9458]  = 211;
  ram[9459]  = 211;
  ram[9460]  = 211;
  ram[9461]  = 211;
  ram[9462]  = 211;
  ram[9463]  = 211;
  ram[9464]  = 211;
  ram[9465]  = 211;
  ram[9466]  = 211;
  ram[9467]  = 211;
  ram[9468]  = 211;
  ram[9469]  = 211;
  ram[9470]  = 211;
  ram[9471]  = 211;
  ram[9472]  = 211;
  ram[9473]  = 211;
  ram[9474]  = 211;
  ram[9475]  = 211;
  ram[9476]  = 211;
  ram[9477]  = 211;
  ram[9478]  = 211;
  ram[9479]  = 211;
  ram[9480]  = 211;
  ram[9481]  = 211;
  ram[9482]  = 211;
  ram[9483]  = 211;
  ram[9484]  = 211;
  ram[9485]  = 211;
  ram[9486]  = 211;
  ram[9487]  = 211;
  ram[9488]  = 211;
  ram[9489]  = 211;
  ram[9490]  = 211;
  ram[9491]  = 211;
  ram[9492]  = 211;
  ram[9493]  = 211;
  ram[9494]  = 211;
  ram[9495]  = 211;
  ram[9496]  = 211;
  ram[9497]  = 211;
  ram[9498]  = 211;
  ram[9499]  = 211;
  ram[9500]  = 211;
  ram[9501]  = 211;
  ram[9502]  = 211;
  ram[9503]  = 211;
  ram[9504]  = 211;
  ram[9505]  = 211;
  ram[9506]  = 211;
  ram[9507]  = 211;
  ram[9508]  = 211;
  ram[9509]  = 211;
  ram[9510]  = 211;
  ram[9511]  = 211;
  ram[9512]  = 211;
  ram[9513]  = 211;
  ram[9514]  = 211;
  ram[9515]  = 211;
  ram[9516]  = 211;
  ram[9517]  = 211;
  ram[9518]  = 211;
  ram[9519]  = 211;
  ram[9520]  = 211;
  ram[9521]  = 211;
  ram[9522]  = 211;
  ram[9523]  = 211;
  ram[9524]  = 211;
  ram[9525]  = 211;
  ram[9526]  = 211;
  ram[9527]  = 211;
  ram[9528]  = 211;
  ram[9529]  = 211;
  ram[9530]  = 211;
  ram[9531]  = 211;
  ram[9532]  = 211;
  ram[9533]  = 211;
  ram[9534]  = 211;
  ram[9535]  = 211;
  ram[9536]  = 211;
  ram[9537]  = 211;
  ram[9538]  = 211;
  ram[9539]  = 211;
  ram[9540]  = 211;
  ram[9541]  = 211;
  ram[9542]  = 211;
  ram[9543]  = 211;
  ram[9544]  = 211;
  ram[9545]  = 211;
  ram[9546]  = 211;
  ram[9547]  = 211;
  ram[9548]  = 211;
  ram[9549]  = 211;
  ram[9550]  = 211;
  ram[9551]  = 211;
  ram[9552]  = 211;
  ram[9553]  = 211;
  ram[9554]  = 211;
  ram[9555]  = 211;
  ram[9556]  = 211;
  ram[9557]  = 211;
  ram[9558]  = 211;
  ram[9559]  = 211;
  ram[9560]  = 211;
  ram[9561]  = 211;
  ram[9562]  = 211;
  ram[9563]  = 211;
  ram[9564]  = 211;
  ram[9565]  = 211;
  ram[9566]  = 211;
  ram[9567]  = 211;
  ram[9568]  = 211;
  ram[9569]  = 211;
  ram[9570]  = 211;
  ram[9571]  = 211;
  ram[9572]  = 211;
  ram[9573]  = 211;
  ram[9574]  = 211;
  ram[9575]  = 211;
  ram[9576]  = 211;
  ram[9577]  = 211;
  ram[9578]  = 211;
  ram[9579]  = 211;
  ram[9580]  = 211;
  ram[9581]  = 211;
  ram[9582]  = 211;
  ram[9583]  = 211;
  ram[9584]  = 211;
  ram[9585]  = 211;
  ram[9586]  = 211;
  ram[9587]  = 211;
  ram[9588]  = 211;
  ram[9589]  = 211;
  ram[9590]  = 211;
  ram[9591]  = 211;
  ram[9592]  = 211;
  ram[9593]  = 210;
  ram[9594]  = 211;
  ram[9595]  = 209;
  ram[9596]  = 208;
  ram[9597]  = 212;
  ram[9598]  = 245;
  ram[9599]  = 255;
  ram[9600]  = 252;
  ram[9601]  = 255;
  ram[9602]  = 255;
  ram[9603]  = 255;
  ram[9604]  = 255;
  ram[9605]  = 255;
  ram[9606]  = 255;
  ram[9607]  = 255;
  ram[9608]  = 255;
  ram[9609]  = 255;
  ram[9610]  = 255;
  ram[9611]  = 255;
  ram[9612]  = 255;
  ram[9613]  = 255;
  ram[9614]  = 255;
  ram[9615]  = 255;
  ram[9616]  = 255;
  ram[9617]  = 255;
  ram[9618]  = 255;
  ram[9619]  = 255;
  ram[9620]  = 255;
  ram[9621]  = 255;
  ram[9622]  = 255;
  ram[9623]  = 255;
  ram[9624]  = 255;
  ram[9625]  = 255;
  ram[9626]  = 255;
  ram[9627]  = 255;
  ram[9628]  = 255;
  ram[9629]  = 255;
  ram[9630]  = 255;
  ram[9631]  = 255;
  ram[9632]  = 255;
  ram[9633]  = 255;
  ram[9634]  = 255;
  ram[9635]  = 255;
  ram[9636]  = 255;
  ram[9637]  = 255;
  ram[9638]  = 255;
  ram[9639]  = 255;
  ram[9640]  = 255;
  ram[9641]  = 255;
  ram[9642]  = 255;
  ram[9643]  = 255;
  ram[9644]  = 255;
  ram[9645]  = 255;
  ram[9646]  = 255;
  ram[9647]  = 255;
  ram[9648]  = 255;
  ram[9649]  = 255;
  ram[9650]  = 255;
  ram[9651]  = 255;
  ram[9652]  = 255;
  ram[9653]  = 255;
  ram[9654]  = 255;
  ram[9655]  = 255;
  ram[9656]  = 255;
  ram[9657]  = 255;
  ram[9658]  = 255;
  ram[9659]  = 255;
  ram[9660]  = 255;
  ram[9661]  = 255;
  ram[9662]  = 255;
  ram[9663]  = 255;
  ram[9664]  = 255;
  ram[9665]  = 255;
  ram[9666]  = 255;
  ram[9667]  = 255;
  ram[9668]  = 255;
  ram[9669]  = 255;
  ram[9670]  = 255;
  ram[9671]  = 255;
  ram[9672]  = 255;
  ram[9673]  = 255;
  ram[9674]  = 255;
  ram[9675]  = 255;
  ram[9676]  = 255;
  ram[9677]  = 255;
  ram[9678]  = 255;
  ram[9679]  = 255;
  ram[9680]  = 255;
  ram[9681]  = 255;
  ram[9682]  = 255;
  ram[9683]  = 255;
  ram[9684]  = 255;
  ram[9685]  = 255;
  ram[9686]  = 255;
  ram[9687]  = 255;
  ram[9688]  = 255;
  ram[9689]  = 255;
  ram[9690]  = 255;
  ram[9691]  = 255;
  ram[9692]  = 255;
  ram[9693]  = 255;
  ram[9694]  = 255;
  ram[9695]  = 255;
  ram[9696]  = 255;
  ram[9697]  = 255;
  ram[9698]  = 255;
  ram[9699]  = 255;
  ram[9700]  = 255;
  ram[9701]  = 255;
  ram[9702]  = 255;
  ram[9703]  = 255;
  ram[9704]  = 255;
  ram[9705]  = 255;
  ram[9706]  = 255;
  ram[9707]  = 255;
  ram[9708]  = 255;
  ram[9709]  = 255;
  ram[9710]  = 255;
  ram[9711]  = 255;
  ram[9712]  = 255;
  ram[9713]  = 255;
  ram[9714]  = 255;
  ram[9715]  = 255;
  ram[9716]  = 255;
  ram[9717]  = 255;
  ram[9718]  = 255;
  ram[9719]  = 255;
  ram[9720]  = 255;
  ram[9721]  = 255;
  ram[9722]  = 255;
  ram[9723]  = 255;
  ram[9724]  = 255;
  ram[9725]  = 255;
  ram[9726]  = 255;
  ram[9727]  = 255;
  ram[9728]  = 255;
  ram[9729]  = 255;
  ram[9730]  = 255;
  ram[9731]  = 255;
  ram[9732]  = 255;
  ram[9733]  = 255;
  ram[9734]  = 255;
  ram[9735]  = 255;
  ram[9736]  = 255;
  ram[9737]  = 255;
  ram[9738]  = 255;
  ram[9739]  = 255;
  ram[9740]  = 255;
  ram[9741]  = 255;
  ram[9742]  = 255;
  ram[9743]  = 255;
  ram[9744]  = 255;
  ram[9745]  = 255;
  ram[9746]  = 255;
  ram[9747]  = 255;
  ram[9748]  = 255;
  ram[9749]  = 255;
  ram[9750]  = 255;
  ram[9751]  = 255;
  ram[9752]  = 255;
  ram[9753]  = 255;
  ram[9754]  = 255;
  ram[9755]  = 255;
  ram[9756]  = 255;
  ram[9757]  = 255;
  ram[9758]  = 255;
  ram[9759]  = 255;
  ram[9760]  = 255;
  ram[9761]  = 255;
  ram[9762]  = 255;
  ram[9763]  = 255;
  ram[9764]  = 255;
  ram[9765]  = 255;
  ram[9766]  = 255;
  ram[9767]  = 255;
  ram[9768]  = 255;
  ram[9769]  = 255;
  ram[9770]  = 255;
  ram[9771]  = 255;
  ram[9772]  = 255;
  ram[9773]  = 255;
  ram[9774]  = 255;
  ram[9775]  = 255;
  ram[9776]  = 255;
  ram[9777]  = 255;
  ram[9778]  = 255;
  ram[9779]  = 255;
  ram[9780]  = 255;
  ram[9781]  = 255;
  ram[9782]  = 255;
  ram[9783]  = 255;
  ram[9784]  = 255;
  ram[9785]  = 255;
  ram[9786]  = 255;
  ram[9787]  = 255;
  ram[9788]  = 255;
  ram[9789]  = 255;
  ram[9790]  = 255;
  ram[9791]  = 255;
  ram[9792]  = 255;
  ram[9793]  = 255;
  ram[9794]  = 255;
  ram[9795]  = 255;
  ram[9796]  = 251;
  ram[9797]  = 255;
  ram[9798]  = 243;
  ram[9799]  = 250;
  ram[9800]  = 249;
  ram[9801]  = 254;
  ram[9802]  = 255;
  ram[9803]  = 255;
  ram[9804]  = 254;
  ram[9805]  = 251;
  ram[9806]  = 247;
  ram[9807]  = 254;
  ram[9808]  = 255;
  ram[9809]  = 255;
  ram[9810]  = 255;
  ram[9811]  = 255;
  ram[9812]  = 255;
  ram[9813]  = 255;
  ram[9814]  = 255;
  ram[9815]  = 255;
  ram[9816]  = 255;
  ram[9817]  = 255;
  ram[9818]  = 255;
  ram[9819]  = 255;
  ram[9820]  = 255;
  ram[9821]  = 255;
  ram[9822]  = 255;
  ram[9823]  = 255;
  ram[9824]  = 255;
  ram[9825]  = 255;
  ram[9826]  = 255;
  ram[9827]  = 255;
  ram[9828]  = 255;
  ram[9829]  = 255;
  ram[9830]  = 255;
  ram[9831]  = 255;
  ram[9832]  = 255;
  ram[9833]  = 255;
  ram[9834]  = 255;
  ram[9835]  = 255;
  ram[9836]  = 255;
  ram[9837]  = 255;
  ram[9838]  = 255;
  ram[9839]  = 255;
  ram[9840]  = 255;
  ram[9841]  = 255;
  ram[9842]  = 255;
  ram[9843]  = 255;
  ram[9844]  = 255;
  ram[9845]  = 255;
  ram[9846]  = 255;
  ram[9847]  = 255;
  ram[9848]  = 255;
  ram[9849]  = 255;
  ram[9850]  = 255;
  ram[9851]  = 255;
  ram[9852]  = 255;
  ram[9853]  = 255;
  ram[9854]  = 255;
  ram[9855]  = 255;
  ram[9856]  = 255;
  ram[9857]  = 255;
  ram[9858]  = 255;
  ram[9859]  = 255;
  ram[9860]  = 255;
  ram[9861]  = 255;
  ram[9862]  = 255;
  ram[9863]  = 255;
  ram[9864]  = 255;
  ram[9865]  = 255;
  ram[9866]  = 255;
  ram[9867]  = 255;
  ram[9868]  = 255;
  ram[9869]  = 255;
  ram[9870]  = 255;
  ram[9871]  = 255;
  ram[9872]  = 255;
  ram[9873]  = 255;
  ram[9874]  = 255;
  ram[9875]  = 255;
  ram[9876]  = 255;
  ram[9877]  = 255;
  ram[9878]  = 255;
  ram[9879]  = 255;
  ram[9880]  = 255;
  ram[9881]  = 255;
  ram[9882]  = 255;
  ram[9883]  = 255;
  ram[9884]  = 255;
  ram[9885]  = 255;
  ram[9886]  = 255;
  ram[9887]  = 255;
  ram[9888]  = 255;
  ram[9889]  = 255;
  ram[9890]  = 255;
  ram[9891]  = 255;
  ram[9892]  = 255;
  ram[9893]  = 255;
  ram[9894]  = 255;
  ram[9895]  = 255;
  ram[9896]  = 255;
  ram[9897]  = 255;
  ram[9898]  = 255;
  ram[9899]  = 255;
  ram[9900]  = 255;
  ram[9901]  = 255;
  ram[9902]  = 255;
  ram[9903]  = 255;
  ram[9904]  = 255;
  ram[9905]  = 255;
  ram[9906]  = 255;
  ram[9907]  = 255;
  ram[9908]  = 255;
  ram[9909]  = 255;
  ram[9910]  = 255;
  ram[9911]  = 255;
  ram[9912]  = 255;
  ram[9913]  = 255;
  ram[9914]  = 255;
  ram[9915]  = 255;
  ram[9916]  = 255;
  ram[9917]  = 255;
  ram[9918]  = 255;
  ram[9919]  = 255;
  ram[9920]  = 255;
  ram[9921]  = 255;
  ram[9922]  = 255;
  ram[9923]  = 255;
  ram[9924]  = 255;
  ram[9925]  = 255;
  ram[9926]  = 255;
  ram[9927]  = 255;
  ram[9928]  = 255;
  ram[9929]  = 255;
  ram[9930]  = 255;
  ram[9931]  = 255;
  ram[9932]  = 255;
  ram[9933]  = 255;
  ram[9934]  = 255;
  ram[9935]  = 255;
  ram[9936]  = 255;
  ram[9937]  = 255;
  ram[9938]  = 255;
  ram[9939]  = 255;
  ram[9940]  = 255;
  ram[9941]  = 255;
  ram[9942]  = 255;
  ram[9943]  = 255;
  ram[9944]  = 255;
  ram[9945]  = 255;
  ram[9946]  = 255;
  ram[9947]  = 255;
  ram[9948]  = 255;
  ram[9949]  = 255;
  ram[9950]  = 255;
  ram[9951]  = 255;
  ram[9952]  = 255;
  ram[9953]  = 255;
  ram[9954]  = 255;
  ram[9955]  = 255;
  ram[9956]  = 255;
  ram[9957]  = 255;
  ram[9958]  = 255;
  ram[9959]  = 255;
  ram[9960]  = 255;
  ram[9961]  = 255;
  ram[9962]  = 255;
  ram[9963]  = 255;
  ram[9964]  = 255;
  ram[9965]  = 255;
  ram[9966]  = 255;
  ram[9967]  = 255;
  ram[9968]  = 255;
  ram[9969]  = 255;
  ram[9970]  = 255;
  ram[9971]  = 255;
  ram[9972]  = 255;
  ram[9973]  = 255;
  ram[9974]  = 255;
  ram[9975]  = 255;
  ram[9976]  = 255;
  ram[9977]  = 255;
  ram[9978]  = 255;
  ram[9979]  = 255;
  ram[9980]  = 255;
  ram[9981]  = 255;
  ram[9982]  = 255;
  ram[9983]  = 255;
  ram[9984]  = 255;
  ram[9985]  = 255;
  ram[9986]  = 255;
  ram[9987]  = 255;
  ram[9988]  = 255;
  ram[9989]  = 255;
  ram[9990]  = 255;
  ram[9991]  = 255;
  ram[9992]  = 255;
  ram[9993]  = 255;
  ram[9994]  = 255;
  ram[9995]  = 255;
  ram[9996]  = 254;
  ram[9997]  = 255;
  ram[9998]  = 253;
  ram[9999]  = 251;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
